// ROM with synchonous read (inferring Block RAM)
// character ROM
//  - 8-by-16 (8-by-2^4) font
//  - 128 (2^7) characters
//  - ROM size: 512-by-8 (2^11-by-8) bits
//              16K bits: 1 BRAM

module font_rom
   (
    input wire clk,
    input wire [12:0] addr,//13 bits
    output reg [31:0] data//32 bits
   );
   
   // signal declaration
   reg [12:0] addr_reg; //13 bits

   // body
   always @(posedge clk) 
      addr_reg <= addr;
      
   always @*
      case (addr_reg)

			//0 x30
						13'h0c00: data = 32'b00000000000000000000000000000000;
						13'h0c01: data = 32'b00000000000011111110000000000000;
						13'h0c02: data = 32'b00000000001111111111100000000000;
						13'h0c03: data = 32'b00000000011111111111110000000000;
						13'h0c04: data = 32'b00000000111111111111111000000000;
						13'h0c05: data = 32'b00000001111111111111111100000000;
						13'h0c06: data = 32'b00000011111111111111111110000000;
						13'h0c07: data = 32'b00000111111111111111111111000000;
						13'h0c08: data = 32'b00000111111111111111111111000000;
						13'h0c09: data = 32'b00001111111111111111111111100000;
						13'h0c0a: data = 32'b00001111111111111111111111100000;
						13'h0c0b: data = 32'b00001111111111111111111111100000;
						13'h0c0c: data = 32'b00011111111110000011111111110000;
						13'h0c0d: data = 32'b00011111111100000001111111110000;
						13'h0c0e: data = 32'b00011111111100000001111111110000;
						13'h0c0f: data = 32'b00111111111000000000111111111000;
						13'h0c10: data = 32'b00111111111000000000111111111000;
						13'h0c11: data = 32'b00111111111000000000111111111000;
						13'h0c12: data = 32'b00111111110000000000011111111000;
						13'h0c13: data = 32'b00111111110000000000011111111000;
						13'h0c14: data = 32'b00111111110000000000011111111000;
						13'h0c15: data = 32'b01111111110000000000011111111100;
						13'h0c16: data = 32'b01111111110000000000011111111100;
						13'h0c17: data = 32'b01111111110000000000011111111100;
						13'h0c18: data = 32'b01111111110000000000011111111100;
						13'h0c19: data = 32'b01111111110000000000011111111100;
						13'h0c1a: data = 32'b01111111110000000000011111111100;
						13'h0c1b: data = 32'b01111111110000000000011111111100;
						13'h0c1c: data = 32'b01111111110000000000011111111100;
						13'h0c1d: data = 32'b01111111110000000000011111111100;
						13'h0c1e: data = 32'b01111111110000000000011111111100;
						13'h0c1f: data = 32'b01111111110000000000011111111100;
						13'h0c20: data = 32'b01111111110000000000011111111100;
						13'h0c21: data = 32'b01111111110000000000011111111100;
						13'h0c22: data = 32'b01111111110000000000011111111100;
						13'h0c23: data = 32'b01111111110000000000011111111100;
						13'h0c24: data = 32'b01111111110000000000011111111100;
						13'h0c25: data = 32'b01111111110000000000011111111100;
						13'h0c26: data = 32'b01111111110000000000011111111100;
						13'h0c27: data = 32'b01111111110000000000011111111100;
						13'h0c28: data = 32'b01111111110000000000011111111100;
						13'h0c29: data = 32'b01111111110000000000011111111100;
						13'h0c2a: data = 32'b00111111110000000000011111111000;
						13'h0c2b: data = 32'b00111111110000000000011111111000;
						13'h0c2c: data = 32'b00111111110000000000011111111000;
						13'h0c2d: data = 32'b00111111111000000000111111111000;
						13'h0c2e: data = 32'b00111111111000000000111111111000;
						13'h0c2f: data = 32'b00111111111000000000111111111000;
						13'h0c30: data = 32'b00011111111000000000111111110000;
						13'h0c31: data = 32'b00011111111100000001111111110000;
						13'h0c32: data = 32'b00011111111100000011111111110000;
						13'h0c33: data = 32'b00011111111111000111111111110000;
						13'h0c34: data = 32'b00001111111111111111111111100000;
						13'h0c35: data = 32'b00001111111111111111111111100000;
						13'h0c36: data = 32'b00000111111111111111111111000000;
						13'h0c37: data = 32'b00000111111111111111111111000000;
						13'h0c38: data = 32'b00000011111111111111111110000000;
						13'h0c39: data = 32'b00000011111111111111111110000000;
						13'h0c3a: data = 32'b00000001111111111111111100000000;
						13'h0c3b: data = 32'b00000000111111111111111000000000;
						13'h0c3c: data = 32'b00000000011111111111110000000000;
						13'h0c3d: data = 32'b00000000000111111111000000000000;
						13'h0c3e: data = 32'b00000000000000111000000000000000;
						13'h0c3f: data = 32'b00000000000000000000000000000000;

			// 1 x32
			13'h0c40: data = 32'b00000000000000000000000000000000;
			13'h0c41: data = 32'b00000000000000000000000000000000;
			13'h0c42: data = 32'b00000000000000001111111110000000;
			13'h0c43: data = 32'b00000000000000001111111110000000;
			13'h0c44: data = 32'b00000000000000011111111110000000;
			13'h0c45: data = 32'b00000000000000011111111110000000;
			13'h0c46: data = 32'b00000000000000111111111110000000;
			13'h0c47: data = 32'b00000000000000111111111110000000;
			13'h0c48: data = 32'b00000000000001111111111110000000;
			13'h0c49: data = 32'b00000000000011111111111110000000;
			13'h0c4a: data = 32'b00000000000111111111111110000000;
			13'h0c4b: data = 32'b00000000001111111111111110000000;
			13'h0c4c: data = 32'b00000000011111111111111110000000;
			13'h0c4d: data = 32'b00000000111111111111111110000000;
			13'h0c4e: data = 32'b00000011111111111111111110000000;
			13'h0c4f: data = 32'b00000111111111111111111110000000;
			13'h0c50: data = 32'b00011111111111111111111110000000;
			13'h0c51: data = 32'b00011111111111111111111110000000;
			13'h0c52: data = 32'b00011111111111111111111110000000;
			13'h0c53: data = 32'b00011111111111011111111110000000;
			13'h0c54: data = 32'b00011111111110011111111110000000;
			13'h0c55: data = 32'b00011111111100011111111110000000;
			13'h0c56: data = 32'b00011111111000011111111110000000;
			13'h0c57: data = 32'b00011111110000011111111110000000;
			13'h0c58: data = 32'b00011111000000011111111110000000;
			13'h0c59: data = 32'b00011100000000011111111110000000;
			13'h0c5a: data = 32'b00010000000000011111111110000000;
			13'h0c5b: data = 32'b00000000000000011111111110000000;
			13'h0c5c: data = 32'b00000000000000011111111110000000;
			13'h0c5d: data = 32'b00000000000000011111111110000000;
			13'h0c5e: data = 32'b00000000000000011111111110000000;
			13'h0c5f: data = 32'b00000000000000011111111110000000;
			13'h0c60: data = 32'b00000000000000011111111110000000;
			13'h0c61: data = 32'b00000000000000011111111110000000;
			13'h0c62: data = 32'b00000000000000011111111110000000;
			13'h0c63: data = 32'b00000000000000011111111110000000;
			13'h0c64: data = 32'b00000000000000011111111110000000;
			13'h0c65: data = 32'b00000000000000011111111110000000;
			13'h0c66: data = 32'b00000000000000011111111110000000;
			13'h0c67: data = 32'b00000000000000011111111110000000;
			13'h0c68: data = 32'b00000000000000011111111110000000;
			13'h0c69: data = 32'b00000000000000011111111110000000;
			13'h0c6a: data = 32'b00000000000000011111111110000000;
			13'h0c6b: data = 32'b00000000000000011111111110000000;
			13'h0c6c: data = 32'b00000000000000011111111110000000;
			13'h0c6d: data = 32'b00000000000000011111111110000000;
			13'h0c6e: data = 32'b00000000000000011111111110000000;
			13'h0c6f: data = 32'b00000000000000011111111110000000;
			13'h0c70: data = 32'b00000000000000011111111110000000;
			13'h0c71: data = 32'b00000000000000011111111110000000;
			13'h0c72: data = 32'b00000000000000011111111110000000;
			13'h0c73: data = 32'b00000000000000011111111110000000;
			13'h0c74: data = 32'b00000000000000011111111110000000;
			13'h0c75: data = 32'b00000000000000011111111110000000;
			13'h0c76: data = 32'b00000000000000011111111110000000;
			13'h0c77: data = 32'b00000000000000011111111110000000;
			13'h0c78: data = 32'b00000000000000011111111110000000;
			13'h0c79: data = 32'b00000000000000011111111110000000;
			13'h0c7a: data = 32'b00000000000000011111111110000000;
			13'h0c7b: data = 32'b00000000000000111111111110000000;
			13'h0c7c: data = 32'b00000000000000000000000000000000;
			13'h0c7d: data = 32'b00000000000000000000000000000000;
			13'h0c7e: data = 32'b00000000000000000000000000000000;
			13'h0c7f: data = 32'b00000000000000000000000000000000;

			//2 x32
			13'h0c80: data = 32'b00000000000000000000000000000000;
			13'h0c81: data = 32'b00000000000000000000000000000000;
			13'h0c82: data = 32'b00000000000000000000000000000000;
			13'h0c83: data = 32'b00000000000011111110000000000000;
			13'h0c84: data = 32'b00000000011111111111111000000000;
			13'h0c85: data = 32'b00000001111111111111111100000000;
			13'h0c86: data = 32'b00000011111111111111111111000000;
			13'h0c87: data = 32'b00000111111111111111111111100000;
			13'h0c88: data = 32'b00001111111111111111111111100000;
			13'h0c89: data = 32'b00011111111111111111111111110000;
			13'h0c8a: data = 32'b00011111111111111111111111111000;
			13'h0c8b: data = 32'b00111111111111111111111111111000;
			13'h0c8c: data = 32'b00111111111111111111111111111000;
			13'h0c8d: data = 32'b00111111111111111111111111111100;
			13'h0c8e: data = 32'b01111111111111111111111111111100;
			13'h0c8f: data = 32'b01111111111111000011111111111100;
			13'h0c90: data = 32'b01111111111110000001111111111100;
			13'h0c91: data = 32'b01111111111100000001111111111110;
			13'h0c92: data = 32'b01111111111100000001111111111110;
			13'h0c93: data = 32'b01111111111100000000111111111110;
			13'h0c94: data = 32'b11111111111100000000111111111110;
			13'h0c95: data = 32'b11111111111000000000111111111110;
			13'h0c96: data = 32'b00001111111000000000111111111110;
			13'h0c97: data = 32'b00000000000000000001111111111100;
			13'h0c98: data = 32'b00000000000000000001111111111100;
			13'h0c99: data = 32'b00000000000000000001111111111100;
			13'h0c9a: data = 32'b00000000000000000011111111111100;
			13'h0c9b: data = 32'b00000000000000000111111111111100;
			13'h0c9c: data = 32'b00000000000000000111111111111000;
			13'h0c9d: data = 32'b00000000000000001111111111111000;
			13'h0c9e: data = 32'b00000000000000011111111111110000;
			13'h0c9f: data = 32'b00000000000000111111111111110000;
			13'h0ca0: data = 32'b00000000000001111111111111100000;
			13'h0ca1: data = 32'b00000000000001111111111111100000;
			13'h0ca2: data = 32'b00000000000011111111111111000000;
			13'h0ca3: data = 32'b00000000000111111111111110000000;
			13'h0ca4: data = 32'b00000000001111111111111110000000;
			13'h0ca5: data = 32'b00000000011111111111111100000000;
			13'h0ca6: data = 32'b00000000111111111111111000000000;
			13'h0ca7: data = 32'b00000000111111111111110000000000;
			13'h0ca8: data = 32'b00000001111111111111100000000000;
			13'h0ca9: data = 32'b00000011111111111111000000000000;
			13'h0caa: data = 32'b00000011111111111110000000000000;
			13'h0cab: data = 32'b00000111111111111110000000000000;
			13'h0cac: data = 32'b00001111111111111100000000000000;
			13'h0cad: data = 32'b00001111111111111000000000000000;
			13'h0cae: data = 32'b00011111111111110000000000000000;
			13'h0caf: data = 32'b00011111111111100000000000000000;
			13'h0cb0: data = 32'b00111111111111111111111111111110;
			13'h0cb1: data = 32'b00111111111111111111111111111110;
			13'h0cb2: data = 32'b00111111111111111111111111111110;
			13'h0cb3: data = 32'b01111111111111111111111111111110;
			13'h0cb4: data = 32'b01111111111111111111111111111110;
			13'h0cb5: data = 32'b01111111111111111111111111111110;
			13'h0cb6: data = 32'b01111111111111111111111111111110;
			13'h0cb7: data = 32'b11111111111111111111111111111110;
			13'h0cb8: data = 32'b11111111111111111111111111111110;
			13'h0cb9: data = 32'b11111111111111111111111111111110;
			13'h0cba: data = 32'b11111111111111111111111111111110;
			13'h0cbb: data = 32'b11111111111111111111111111111110;
			13'h0cbc: data = 32'b11111111111111111111111111111110;
			13'h0cbd: data = 32'b00000000000000000000000000000000;
			13'h0cbe: data = 32'b00000000000000000000000000000000;
			13'h0cbf: data = 32'b00000000000000000000000000000000;

			//3 x33
			13'h0cc0: data = 32'b00000000000000000000000000000000;
			13'h0cc1: data = 32'b00000000000000111100000000000000;
			13'h0cc2: data = 32'b00000000000111111111100000000000;
			13'h0cc3: data = 32'b00000000001111111111110000000000;
			13'h0cc4: data = 32'b00000000011111111111111000000000;
			13'h0cc5: data = 32'b00000000111111111111111100000000;
			13'h0cc6: data = 32'b00000001111111111111111110000000;
			13'h0cc7: data = 32'b00000011111111111111111110000000;
			13'h0cc8: data = 32'b00000011111111111111111111000000;
			13'h0cc9: data = 32'b00000111111111111111111111000000;
			13'h0cca: data = 32'b00000111111111111111111111100000;
			13'h0ccb: data = 32'b00000111111111100111111111100000;
			13'h0ccc: data = 32'b00000111111110000011111111100000;
			13'h0ccd: data = 32'b00001111111110000001111111100000;
			13'h0cce: data = 32'b00001111111100000001111111100000;
			13'h0ccf: data = 32'b00001111111100000001111111110000;
			13'h0cd0: data = 32'b00001111111100000001111111110000;
			13'h0cd1: data = 32'b00000111111000000001111111110000;
			13'h0cd2: data = 32'b00000000111000000001111111110000;
			13'h0cd3: data = 32'b00000000000000000001111111100000;
			13'h0cd4: data = 32'b00000000000000000001111111100000;
			13'h0cd5: data = 32'b00000000000000000001111111100000;
			13'h0cd6: data = 32'b00000000000000000011111111100000;
			13'h0cd7: data = 32'b00000000000000000111111111000000;
			13'h0cd8: data = 32'b00000000000000011111111111000000;
			13'h0cd9: data = 32'b00000000000001111111111110000000;
			13'h0cda: data = 32'b00000000000001111111111110000000;
			13'h0cdb: data = 32'b00000000000001111111111100000000;
			13'h0cdc: data = 32'b00000000000001111111111000000000;
			13'h0cdd: data = 32'b00000000000001111111111100000000;
			13'h0cde: data = 32'b00000000000001111111111110000000;
			13'h0cdf: data = 32'b00000000000001111111111111000000;
			13'h0ce0: data = 32'b00000000000001111111111111100000;
			13'h0ce1: data = 32'b00000000000001111111111111100000;
			13'h0ce2: data = 32'b00000000000000000001111111110000;
			13'h0ce3: data = 32'b00000000000000000000111111110000;
			13'h0ce4: data = 32'b00000000000000000000111111110000;
			13'h0ce5: data = 32'b00000000000000000000111111111000;
			13'h0ce6: data = 32'b00000000000000000000011111111000;
			13'h0ce7: data = 32'b00000000000000000000011111111000;
			13'h0ce8: data = 32'b00000000000000000000011111111000;
			13'h0ce9: data = 32'b00000000000000000000011111111000;
			13'h0cea: data = 32'b00000000000000000000011111111000;
			13'h0ceb: data = 32'b00000000111000000000011111111000;
			13'h0cec: data = 32'b00011111111000000000011111111000;
			13'h0ced: data = 32'b00011111111000000000011111111000;
			13'h0cee: data = 32'b00011111111100000000011111111000;
			13'h0cef: data = 32'b00001111111100000000111111111000;
			13'h0cf0: data = 32'b00001111111100000000111111111000;
			13'h0cf1: data = 32'b00001111111110000001111111111000;
			13'h0cf2: data = 32'b00001111111110000001111111110000;
			13'h0cf3: data = 32'b00000111111111100111111111110000;
			13'h0cf4: data = 32'b00000111111111111111111111100000;
			13'h0cf5: data = 32'b00000111111111111111111111100000;
			13'h0cf6: data = 32'b00000011111111111111111111100000;
			13'h0cf7: data = 32'b00000011111111111111111111000000;
			13'h0cf8: data = 32'b00000001111111111111111110000000;
			13'h0cf9: data = 32'b00000000111111111111111100000000;
			13'h0cfa: data = 32'b00000000011111111111111100000000;
			13'h0cfb: data = 32'b00000000001111111111110000000000;
			13'h0cfc: data = 32'b00000000000111111111100000000000;
			13'h0cfd: data = 32'b00000000000000111100000000000000;
			13'h0cfe: data = 32'b00000000000000000000000000000000;
			13'h0cff: data = 32'b00000000000000000000000000000000;

			//4 x34
			13'h0d00: data = 32'b00000000000000000000000000000000;
			13'h0d01: data = 32'b00000000000000000000000000000000;
			13'h0d02: data = 32'b00000000000000000000000000000000;
			13'h0d03: data = 32'b00000000000000000000000000000000;
			13'h0d04: data = 32'b00000000000000000000000000000000;
			13'h0d05: data = 32'b00000000000000000000000000000000;
			13'h0d06: data = 32'b00000000000000000000000000000000;
			13'h0d07: data = 32'b00000000000000000000000000000000;
			13'h0d08: data = 32'b00000000000000000001111110000000;
			13'h0d09: data = 32'b00000000000000000001111110000000;
			13'h0d0a: data = 32'b00000000000000000001111110000000;
			13'h0d0b: data = 32'b00000000000000000011111110000000;
			13'h0d0c: data = 32'b00000000000000000011111110000000;
			13'h0d0d: data = 32'b00000000000000000111111110000000;
			13'h0d0e: data = 32'b00000000000000000111111110000000;
			13'h0d0f: data = 32'b00000000000000001111111110000000;
			13'h0d10: data = 32'b00000000000000001111111110000000;
			13'h0d11: data = 32'b00000000000000001111111110000000;
			13'h0d12: data = 32'b00000000000000011111111110000000;
			13'h0d13: data = 32'b00000000000000011111111110000000;
			13'h0d14: data = 32'b00000000000000111111111110000000;
			13'h0d15: data = 32'b00000000000000111111111110000000;
			13'h0d16: data = 32'b00000000000001111110111110000000;
			13'h0d17: data = 32'b00000000000001111110111110000000;
			13'h0d18: data = 32'b00000000000001111100111110000000;
			13'h0d19: data = 32'b00000000000011111100111110000000;
			13'h0d1a: data = 32'b00000000000011111100111110000000;
			13'h0d1b: data = 32'b00000000000111111000111110000000;
			13'h0d1c: data = 32'b00000000000111111000111110000000;
			13'h0d1d: data = 32'b00000000001111110000111110000000;
			13'h0d1e: data = 32'b00000000001111110000111110000000;
			13'h0d1f: data = 32'b00000000001111100000111110000000;
			13'h0d20: data = 32'b00000000011111100000111110000000;
			13'h0d21: data = 32'b00000000011111100000111110000000;
			13'h0d22: data = 32'b00000000111111000000111110000000;
			13'h0d23: data = 32'b00000000111111000000111110000000;
			13'h0d24: data = 32'b00000000111110000000111110000000;
			13'h0d25: data = 32'b00000001111110000000111110000000;
			13'h0d26: data = 32'b00000001111100000000111110000000;
			13'h0d27: data = 32'b00000011111111111111111111110000;
			13'h0d28: data = 32'b00000011111111111111111111110000;
			13'h0d29: data = 32'b00000111111111111111111111110000;
			13'h0d2a: data = 32'b00000111111111111111111111110000;
			13'h0d2b: data = 32'b00000111111111111111111111110000;
			13'h0d2c: data = 32'b00000111111111111111111111110000;
			13'h0d2d: data = 32'b00000111111111111111111111110000;
			13'h0d2e: data = 32'b00000111111111111111111111110000;
			13'h0d2f: data = 32'b00000000000000000000111110000000;
			13'h0d30: data = 32'b00000000000000000000111110000000;
			13'h0d31: data = 32'b00000000000000000000111110000000;
			13'h0d32: data = 32'b00000000000000000000111110000000;
			13'h0d33: data = 32'b00000000000000000000111110000000;
			13'h0d34: data = 32'b00000000000000000000111110000000;
			13'h0d35: data = 32'b00000000000000000000111110000000;
			13'h0d36: data = 32'b00000000000000000000111110000000;
			13'h0d37: data = 32'b00000000000000000000111110000000;
			13'h0d38: data = 32'b00000000000000000000111110000000;
			13'h0d39: data = 32'b00000000000000000000111110000000;
			13'h0d3a: data = 32'b00000000000000000000111110000000;
			13'h0d3b: data = 32'b00000000000000000000111110000000;
			13'h0d3c: data = 32'b00000000000000000000000000000000;
			13'h0d3d: data = 32'b00000000000000000000000000000000;
			13'h0d3e: data = 32'b00000000000000000000000000000000;
			13'h0d3f: data = 32'b00000000000000000000000000000000;

			//5 x35
			13'h0d40: data = 32'b00000000000000000000000000000000;
			13'h0d41: data = 32'b00000000000000000000000000000000;
			13'h0d42: data = 32'b00000000000000000000000000000000;
			13'h0d43: data = 32'b00000000000000000000000000000000;
			13'h0d44: data = 32'b00000011111111111111111111000000;
			13'h0d45: data = 32'b00000011111111111111111111000000;
			13'h0d46: data = 32'b00000011111111111111111111000000;
			13'h0d47: data = 32'b00000011111111111111111111000000;
			13'h0d48: data = 32'b00000011111111111111111111000000;
			13'h0d49: data = 32'b00000011111111111111111111000000;
			13'h0d4a: data = 32'b00000111111111111111111111000000;
			13'h0d4b: data = 32'b00000111111111111111111111000000;
			13'h0d4c: data = 32'b00000111111111111111111111000000;
			13'h0d4d: data = 32'b00000111111111111111111111000000;
			13'h0d4e: data = 32'b00000111111111111111111111000000;
			13'h0d4f: data = 32'b00000111111100000000000000000000;
			13'h0d50: data = 32'b00000111111100000000000000000000;
			13'h0d51: data = 32'b00000111111100000000000000000000;
			13'h0d52: data = 32'b00001111111100000000000000000000;
			13'h0d53: data = 32'b00001111111100000000000000000000;
			13'h0d54: data = 32'b00001111111100000000000000000000;
			13'h0d55: data = 32'b00001111111100000000000000000000;
			13'h0d56: data = 32'b00001111111101111111000000000000;
			13'h0d57: data = 32'b00001111111111111111100000000000;
			13'h0d58: data = 32'b00001111111111111111111000000000;
			13'h0d59: data = 32'b00001111111111111111111100000000;
			13'h0d5a: data = 32'b00011111111111111111111100000000;
			13'h0d5b: data = 32'b00011111111111111111111110000000;
			13'h0d5c: data = 32'b00011111111111111111111111000000;
			13'h0d5d: data = 32'b00011111111111111111111111000000;
			13'h0d5e: data = 32'b00011111111111111111111111000000;
			13'h0d5f: data = 32'b00011111111100000111111111100000;
			13'h0d60: data = 32'b00011111111000000011111111100000;
			13'h0d61: data = 32'b00011111110000000011111111100000;
			13'h0d62: data = 32'b00000011100000000001111111110000;
			13'h0d63: data = 32'b00000000000000000001111111110000;
			13'h0d64: data = 32'b00000000000000000001111111110000;
			13'h0d65: data = 32'b00000000000000000000111111110000;
			13'h0d66: data = 32'b00000000000000000000111111110000;
			13'h0d67: data = 32'b00000000000000000000111111110000;
			13'h0d68: data = 32'b00000000000000000000111111110000;
			13'h0d69: data = 32'b00000000000000000000111111110000;
			13'h0d6a: data = 32'b00000000000000000000111111110000;
			13'h0d6b: data = 32'b00000000000000000000111111110000;
			13'h0d6c: data = 32'b00000111110000000000111111110000;
			13'h0d6d: data = 32'b00111111110000000000111111110000;
			13'h0d6e: data = 32'b00111111110000000001111111110000;
			13'h0d6f: data = 32'b00111111110000000001111111100000;
			13'h0d70: data = 32'b00111111111000000001111111100000;
			13'h0d71: data = 32'b00111111111000000011111111100000;
			13'h0d72: data = 32'b00011111111100000011111111100000;
			13'h0d73: data = 32'b00011111111110001111111111000000;
			13'h0d74: data = 32'b00011111111111111111111111000000;
			13'h0d75: data = 32'b00001111111111111111111110000000;
			13'h0d76: data = 32'b00001111111111111111111110000000;
			13'h0d77: data = 32'b00000111111111111111111100000000;
			13'h0d78: data = 32'b00000111111111111111111100000000;
			13'h0d79: data = 32'b00000011111111111111111000000000;
			13'h0d7a: data = 32'b00000001111111111111110000000000;
			13'h0d7b: data = 32'b00000000011111111111100000000000;
			13'h0d7c: data = 32'b00000000001111111110000000000000;
			13'h0d7d: data = 32'b00000000000000000000000000000000;
			13'h0d7e: data = 32'b00000000000000000000000000000000;
			13'h0d7f: data = 32'b00000000000000000000000000000000;

			//6 x36
			13'h0d80: data = 32'b00000000000000000000000000000000;
			13'h0d81: data = 32'b00000000000001111100000000000000;
			13'h0d82: data = 32'b00000000000111111111000000000000;
			13'h0d83: data = 32'b00000000011111111111100000000000;
			13'h0d84: data = 32'b00000000111111111111110000000000;
			13'h0d85: data = 32'b00000000111111111111111000000000;
			13'h0d86: data = 32'b00000001111111111111111100000000;
			13'h0d87: data = 32'b00000011111111111111111100000000;
			13'h0d88: data = 32'b00000011111111111111111110000000;
			13'h0d89: data = 32'b00000111111111111111111110000000;
			13'h0d8a: data = 32'b00000111111111111111111110000000;
			13'h0d8b: data = 32'b00001111111111001111111111000000;
			13'h0d8c: data = 32'b00001111111110000111111111000000;
			13'h0d8d: data = 32'b00001111111100000011111111000000;
			13'h0d8e: data = 32'b00011111111100000011111111000000;
			13'h0d8f: data = 32'b00011111111000000001111111000000;
			13'h0d90: data = 32'b00011111111000000001111111000000;
			13'h0d91: data = 32'b00011111111000000001100000000000;
			13'h0d92: data = 32'b00011111111000000000000000000000;
			13'h0d93: data = 32'b00111111110000000000000000000000;
			13'h0d94: data = 32'b00111111110000000000000000000000;
			13'h0d95: data = 32'b00111111110000000000000000000000;
			13'h0d96: data = 32'b00111111110001111110000000000000;
			13'h0d97: data = 32'b00111111110011111111000000000000;
			13'h0d98: data = 32'b00111111110111111111110000000000;
			13'h0d99: data = 32'b00111111111111111111110000000000;
			13'h0d9a: data = 32'b00111111111111111111111000000000;
			13'h0d9b: data = 32'b00111111111111111111111100000000;
			13'h0d9c: data = 32'b00111111111111111111111100000000;
			13'h0d9d: data = 32'b00111111111111111111111110000000;
			13'h0d9e: data = 32'b00111111111111111111111110000000;
			13'h0d9f: data = 32'b00111111111110000111111111000000;
			13'h0da0: data = 32'b00111111111100000011111111000000;
			13'h0da1: data = 32'b00111111111100000011111111000000;
			13'h0da2: data = 32'b00111111111000000001111111000000;
			13'h0da3: data = 32'b00111111111000000001111111100000;
			13'h0da4: data = 32'b00111111111000000001111111100000;
			13'h0da5: data = 32'b00111111111000000001111111100000;
			13'h0da6: data = 32'b00111111110000000001111111100000;
			13'h0da7: data = 32'b00111111110000000001111111100000;
			13'h0da8: data = 32'b00111111110000000001111111100000;
			13'h0da9: data = 32'b00111111110000000001111111100000;
			13'h0daa: data = 32'b00111111110000000001111111100000;
			13'h0dab: data = 32'b00111111111000000001111111100000;
			13'h0dac: data = 32'b00011111111000000001111111100000;
			13'h0dad: data = 32'b00011111111000000001111111100000;
			13'h0dae: data = 32'b00011111111000000001111111100000;
			13'h0daf: data = 32'b00011111111000000001111111100000;
			13'h0db0: data = 32'b00011111111100000011111111000000;
			13'h0db1: data = 32'b00001111111100000011111111000000;
			13'h0db2: data = 32'b00001111111110000111111111000000;
			13'h0db3: data = 32'b00001111111111111111111111000000;
			13'h0db4: data = 32'b00000111111111111111111110000000;
			13'h0db5: data = 32'b00000111111111111111111110000000;
			13'h0db6: data = 32'b00000111111111111111111100000000;
			13'h0db7: data = 32'b00000011111111111111111100000000;
			13'h0db8: data = 32'b00000001111111111111111000000000;
			13'h0db9: data = 32'b00000001111111111111110000000000;
			13'h0dba: data = 32'b00000000111111111111110000000000;
			13'h0dbb: data = 32'b00000000011111111111000000000000;
			13'h0dbc: data = 32'b00000000000111111110000000000000;
			13'h0dbd: data = 32'b00000000000000000000000000000000;
			13'h0dbe: data = 32'b00000000000000000000000000000000;
			13'h0dbf: data = 32'b00000000000000000000000000000000;

			// 7 x37
			13'h0dc0: data = 32'b00000000000000000000000000000000;
			13'h0dc1: data = 32'b00111111111111111111111111111000;
			13'h0dc2: data = 32'b00111111111111111111111111111000;
			13'h0dc3: data = 32'b00111111111111111111111111111000;
			13'h0dc4: data = 32'b00111111111111111111111111111000;
			13'h0dc5: data = 32'b00111111111111111111111111111000;
			13'h0dc6: data = 32'b00111111111111111111111111111000;
			13'h0dc7: data = 32'b00111111111111111111111111111000;
			13'h0dc8: data = 32'b00111111111111111111111111111000;
			13'h0dc9: data = 32'b00111111111111111111111111111000;
			13'h0dca: data = 32'b00111111111111111111111111111000;
			13'h0dcb: data = 32'b00111111111111111111111111111000;
			13'h0dcc: data = 32'b00111111111111111111111111111000;
			13'h0dcd: data = 32'b00111111111111111111111111111000;
			13'h0dce: data = 32'b00111111111111111111111111111000;
			13'h0dcf: data = 32'b00111111111000000011111111111000;
			13'h0dd0: data = 32'b00111111111000000011111111111000;
			13'h0dd1: data = 32'b00111111111000000111111111110000;
			13'h0dd2: data = 32'b00111111111000000111111111110000;
			13'h0dd3: data = 32'b00000000000000000111111111110000;
			13'h0dd4: data = 32'b00000000000000000111111111110000;
			13'h0dd5: data = 32'b00000000000000001111111111100000;
			13'h0dd6: data = 32'b00000000000000001111111111100000;
			13'h0dd7: data = 32'b00000000000000001111111111100000;
			13'h0dd8: data = 32'b00000000000000001111111111100000;
			13'h0dd9: data = 32'b00000000000000001111111111100000;
			13'h0dda: data = 32'b00000000000000011111111111000000;
			13'h0ddb: data = 32'b00000000000000011111111111000000;
			13'h0ddc: data = 32'b00000000000000011111111111000000;
			13'h0ddd: data = 32'b00000000000000011111111111000000;
			13'h0dde: data = 32'b00000000000000011111111111000000;
			13'h0ddf: data = 32'b00000000000000111111111110000000;
			13'h0de0: data = 32'b00000000000000111111111110000000;
			13'h0de1: data = 32'b00000000000000111111111110000000;
			13'h0de2: data = 32'b00000000000000111111111110000000;
			13'h0de3: data = 32'b00000000000001111111111100000000;
			13'h0de4: data = 32'b00000000000001111111111100000000;
			13'h0de5: data = 32'b00000000000001111111111100000000;
			13'h0de6: data = 32'b00000000000001111111111100000000;
			13'h0de7: data = 32'b00000000000001111111111100000000;
			13'h0de8: data = 32'b00000000000011111111111000000000;
			13'h0de9: data = 32'b00000000000011111111111000000000;
			13'h0dea: data = 32'b00000000000011111111111000000000;
			13'h0deb: data = 32'b00000000000011111111111000000000;
			13'h0dec: data = 32'b00000000000111111111110000000000;
			13'h0ded: data = 32'b00000000000111111111110000000000;
			13'h0dee: data = 32'b00000000000111111111110000000000;
			13'h0def: data = 32'b00000000000111111111110000000000;
			13'h0df0: data = 32'b00000000000111111111110000000000;
			13'h0df1: data = 32'b00000000001111111111100000000000;
			13'h0df2: data = 32'b00000000001111111111100000000000;
			13'h0df3: data = 32'b00000000001111111111100000000000;
			13'h0df4: data = 32'b00000000001111111111100000000000;
			13'h0df5: data = 32'b00000000001111111111000000000000;
			13'h0df6: data = 32'b00000000011111111111000000000000;
			13'h0df7: data = 32'b00000000011111111111000000000000;
			13'h0df8: data = 32'b00000000011111111111000000000000;
			13'h0df9: data = 32'b00000000011111111111000000000000;
			13'h0dfa: data = 32'b00000000111111111110000000000000;
			13'h0dfb: data = 32'b00000000111111111110000000000000;
			13'h0dfc: data = 32'b00000000111111111110000000000000;
			13'h0dfd: data = 32'b00000000111111111110000000000000;
			13'h0dfe: data = 32'b00000000111111111110000000000000;
			13'h0dff: data = 32'b00000000000000000000000000000000;

			// 8 x38
			13'h0e00: data = 32'b00000000000000000000000000000000;
			13'h0e01: data = 32'b00000000000111111110000000000000;
			13'h0e02: data = 32'b00000000011111111111000000000000;
			13'h0e03: data = 32'b00000000111111111111100000000000;
			13'h0e04: data = 32'b00000001111111111111110000000000;
			13'h0e05: data = 32'b00000001111111111111111000000000;
			13'h0e06: data = 32'b00000011111111111111111000000000;
			13'h0e07: data = 32'b00000011111111111111111100000000;
			13'h0e08: data = 32'b00000111111111111111111100000000;
			13'h0e09: data = 32'b00000111111111111111111100000000;
			13'h0e0a: data = 32'b00000111111111111111111110000000;
			13'h0e0b: data = 32'b00000111111110000111111110000000;
			13'h0e0c: data = 32'b00001111111100000011111110000000;
			13'h0e0d: data = 32'b00001111111100000011111110000000;
			13'h0e0e: data = 32'b00001111111000000011111110000000;
			13'h0e0f: data = 32'b00001111111000000011111110000000;
			13'h0e10: data = 32'b00001111111000000011111110000000;
			13'h0e11: data = 32'b00001111111000000011111110000000;
			13'h0e12: data = 32'b00001111111000000011111110000000;
			13'h0e13: data = 32'b00001111111000000011111110000000;
			13'h0e14: data = 32'b00000111111000000011111110000000;
			13'h0e15: data = 32'b00000111111100000011111110000000;
			13'h0e16: data = 32'b00000111111100000111111110000000;
			13'h0e17: data = 32'b00000111111110000111111100000000;
			13'h0e18: data = 32'b00000011111111111111111100000000;
			13'h0e19: data = 32'b00000011111111111111111000000000;
			13'h0e1a: data = 32'b00000001111111111111111000000000;
			13'h0e1b: data = 32'b00000001111111111111110000000000;
			13'h0e1c: data = 32'b00000000011111111111100000000000;
			13'h0e1d: data = 32'b00000000111111111111110000000000;
			13'h0e1e: data = 32'b00000001111111111111111000000000;
			13'h0e1f: data = 32'b00000011111111111111111000000000;
			13'h0e20: data = 32'b00000011111111111111111100000000;
			13'h0e21: data = 32'b00000111111111111111111100000000;
			13'h0e22: data = 32'b00000111111110001111111110000000;
			13'h0e23: data = 32'b00000111111100000111111110000000;
			13'h0e24: data = 32'b00001111111100000011111111000000;
			13'h0e25: data = 32'b00001111111000000011111111000000;
			13'h0e26: data = 32'b00001111111000000001111111000000;
			13'h0e27: data = 32'b00001111111000000001111111000000;
			13'h0e28: data = 32'b00001111111000000001111111000000;
			13'h0e29: data = 32'b00011111111000000001111111000000;
			13'h0e2a: data = 32'b00011111111000000001111111000000;
			13'h0e2b: data = 32'b00011111111000000001111111000000;
			13'h0e2c: data = 32'b00011111111000000001111111000000;
			13'h0e2d: data = 32'b00011111111000000001111111000000;
			13'h0e2e: data = 32'b00011111111000000001111111000000;
			13'h0e2f: data = 32'b00011111111000000001111111000000;
			13'h0e30: data = 32'b00001111111000000001111111000000;
			13'h0e31: data = 32'b00001111111000000011111111000000;
			13'h0e32: data = 32'b00001111111100000011111111000000;
			13'h0e33: data = 32'b00001111111110000111111111000000;
			13'h0e34: data = 32'b00001111111111001111111110000000;
			13'h0e35: data = 32'b00000111111111111111111110000000;
			13'h0e36: data = 32'b00000111111111111111111110000000;
			13'h0e37: data = 32'b00000011111111111111111100000000;
			13'h0e38: data = 32'b00000011111111111111111100000000;
			13'h0e39: data = 32'b00000001111111111111111000000000;
			13'h0e3a: data = 32'b00000001111111111111111000000000;
			13'h0e3b: data = 32'b00000000111111111111110000000000;
			13'h0e3c: data = 32'b00000000011111111111100000000000;
			13'h0e3d: data = 32'b00000000000111111110000000000000;
			13'h0e3e: data = 32'b00000000000001111000000000000000;
			13'h0e3f: data = 32'b00000000000000000000000000000000;

			// 9 x39
			13'h0e40: data = 32'b00000000000000000000000000000000;
			13'h0e41: data = 32'b00000000000000000000000000000000;
			13'h0e42: data = 32'b00000000000000110000000000000000;
			13'h0e43: data = 32'b00000000000111111110000000000000;
			13'h0e44: data = 32'b00000000001111111111000000000000;
			13'h0e45: data = 32'b00000000011111111111100000000000;
			13'h0e46: data = 32'b00000000111111111111110000000000;
			13'h0e47: data = 32'b00000001111111111111111000000000;
			13'h0e48: data = 32'b00000001111111111111111000000000;
			13'h0e49: data = 32'b00000011111111111111111100000000;
			13'h0e4a: data = 32'b00000011111111111111111100000000;
			13'h0e4b: data = 32'b00000111111111111111111110000000;
			13'h0e4c: data = 32'b00000111111111001111111110000000;
			13'h0e4d: data = 32'b00000111111110000111111110000000;
			13'h0e4e: data = 32'b00001111111100000011111111000000;
			13'h0e4f: data = 32'b00001111111100000011111111000000;
			13'h0e50: data = 32'b00001111111000000011111111000000;
			13'h0e51: data = 32'b00001111111000000001111111000000;
			13'h0e52: data = 32'b00001111111000000001111111000000;
			13'h0e53: data = 32'b00001111111000000001111111100000;
			13'h0e54: data = 32'b00001111111000000001111111100000;
			13'h0e55: data = 32'b00001111111000000001111111100000;
			13'h0e56: data = 32'b00001111111000000001111111100000;
			13'h0e57: data = 32'b00001111111000000001111111100000;
			13'h0e58: data = 32'b00001111111000000001111111100000;
			13'h0e59: data = 32'b00001111111000000001111111100000;
			13'h0e5a: data = 32'b00001111111000000001111111100000;
			13'h0e5b: data = 32'b00001111111000000001111111100000;
			13'h0e5c: data = 32'b00001111111100000001111111100000;
			13'h0e5d: data = 32'b00000111111100000011111111100000;
			13'h0e5e: data = 32'b00000111111110000011111111100000;
			13'h0e5f: data = 32'b00000111111110000111111111100000;
			13'h0e60: data = 32'b00000111111111111111111111100000;
			13'h0e61: data = 32'b00000011111111111111111111100000;
			13'h0e62: data = 32'b00000011111111111111111111100000;
			13'h0e63: data = 32'b00000001111111111111111111100000;
			13'h0e64: data = 32'b00000001111111111111111111100000;
			13'h0e65: data = 32'b00000000111111111110111111100000;
			13'h0e66: data = 32'b00000000011111111110111111100000;
			13'h0e67: data = 32'b00000000001111111100111111100000;
			13'h0e68: data = 32'b00000000000011110001111111100000;
			13'h0e69: data = 32'b00000000000000000001111111100000;
			13'h0e6a: data = 32'b00000000000000000001111111100000;
			13'h0e6b: data = 32'b00000000000000000001111111100000;
			13'h0e6c: data = 32'b00000000000000000001111111000000;
			13'h0e6d: data = 32'b00000000111100000001111111000000;
			13'h0e6e: data = 32'b00001111111100000001111111000000;
			13'h0e6f: data = 32'b00000111111100000011111111000000;
			13'h0e70: data = 32'b00000111111100000011111111000000;
			13'h0e71: data = 32'b00000111111100000111111110000000;
			13'h0e72: data = 32'b00000111111110000111111110000000;
			13'h0e73: data = 32'b00000111111111111111111110000000;
			13'h0e74: data = 32'b00000011111111111111111100000000;
			13'h0e75: data = 32'b00000011111111111111111100000000;
			13'h0e76: data = 32'b00000011111111111111111000000000;
			13'h0e77: data = 32'b00000001111111111111111000000000;
			13'h0e78: data = 32'b00000001111111111111110000000000;
			13'h0e79: data = 32'b00000000111111111111100000000000;
			13'h0e7a: data = 32'b00000000011111111111000000000000;
			13'h0e7b: data = 32'b00000000001111111110000000000000;
			13'h0e7c: data = 32'b00000000000011111000000000000000;
			13'h0e7d: data = 32'b00000000000000000000000000000000;
			13'h0e7e: data = 32'b00000000000000000000000000000000;
			13'h0e7f: data = 32'b00000000000000000000000000000000;

		
// A x40
         13'h1040: data = 32'b00000000000000000000000000000000;
			13'h1041: data = 32'b00000000000000000000000000000000;
			13'h1042: data = 32'b00000000000000000000000000000000;
			13'h1043: data = 32'b00000000000000000000000000000000;
			13'h1044: data = 32'b00000000000000000000000000000000;
			13'h1045: data = 32'b00000000000000000000000000000000;
			13'h1046: data = 32'b00000000000000000000000000000000;
			13'h1047: data = 32'b00000000000000000000000000000000;
			13'h1048: data = 32'b00000000000001111111000000000000;
			13'h1049: data = 32'b00000000000001111111000000000000;
			13'h104a: data = 32'b00000000000011111111000000000000;
			13'h104b: data = 32'b00000000000111111111100000000000;
			13'h104c: data = 32'b00000000000111111111100000000000;
			13'h104d: data = 32'b00000000000111111111100000000000;
			13'h104e: data = 32'b00000000000111111111100000000000;
			13'h104f: data = 32'b00000000000111111111100000000000;
			13'h1050: data = 32'b00000000001111111111110000000000;
			13'h1051: data = 32'b00000000001111111111110000000000;
			13'h1052: data = 32'b00000000001111111111110000000000;
			13'h1053: data = 32'b00000000001111111111110000000000;
			13'h1054: data = 32'b00000000011111111111111000000000;
			13'h1055: data = 32'b00000000011111111111111000000000;
			13'h1056: data = 32'b00000000011111111111111000000000;
			13'h1057: data = 32'b00000000011111111111111000000000;
			13'h1058: data = 32'b00000000011111111111111000000000;
			13'h1059: data = 32'b00000000011111111111111100000000;
			13'h105a: data = 32'b00000000011111111111111100000000;
			13'h105b: data = 32'b00000000011111111111111100000000;
			13'h105c: data = 32'b00000000111111111111111110000000;
			13'h105d: data = 32'b00000000111111111111111110000000;
			13'h105e: data = 32'b00000000111111100111111110000000;
			13'h105f: data = 32'b00000000111111100111111110000000;
			13'h1060: data = 32'b00000000111111100111111110000000;
			13'h1061: data = 32'b00000000111111100111111110000000;
			13'h1062: data = 32'b00000001111111100111111111000000;
			13'h1063: data = 32'b00000001111111000011111111000000;
			13'h1064: data = 32'b00000001111111000011111111000000;
			13'h1065: data = 32'b00000001111111000011111111000000;
			13'h1066: data = 32'b00000001111111000011111111000000;
			13'h1067: data = 32'b00000011111111000011111111100000;
			13'h1068: data = 32'b00000111111111111111111111100000;
			13'h1069: data = 32'b00000111111111111111111111100000;
			13'h106a: data = 32'b00000111111111111111111111100000;
			13'h106b: data = 32'b00000111111111111111111111100000;
			13'h106c: data = 32'b00000111111111111111111111100000;
			13'h106d: data = 32'b00001111111111111111111111110000;
			13'h106e: data = 32'b00001111111111111111111111110000;
			13'h106f: data = 32'b00001111111111111111111111110000;
			13'h1070: data = 32'b00001111111111111111111111110000;
			13'h1071: data = 32'b00001111111111111111111111110000;
			13'h1072: data = 32'b00011111111111111111111111111000;
			13'h1073: data = 32'b00011111111100000000111111111000;
			13'h1074: data = 32'b00011111111000000000011111111000;
			13'h1075: data = 32'b00011111111000000000011111111000;
			13'h1076: data = 32'b00011111111000000000011111111000;
			13'h1077: data = 32'b00111111111000000000011111111100;
			13'h1078: data = 32'b00111111111000000000011111111100;
			13'h1079: data = 32'b00111111111000000000011111111100;
			13'h107a: data = 32'b00111111111000000000011111111100;
			13'h107b: data = 32'b00000000000000000000000000000000;
			13'h107c: data = 32'b00000000000000000000000000000000;
			13'h107d: data = 32'b00000000000000000000000000000000;
			13'h107e: data = 32'b00000000000000000000000000000000;
			13'h107f: data = 32'b00000000000000000000000000000000; 
         
//B x42
			13'h1080: data = 32'b00000000000000000000000000000000;
			13'h1081: data = 32'b00000000000000000000000000000000;
			13'h1082: data = 32'b00000000000000000000000000000000;
			13'h1083: data = 32'b00000000000000000000000000000000;
			13'h1084: data = 32'b00000000000000000000000000000000;
			13'h1085: data = 32'b00000000000000000000000000000000;
			13'h1086: data = 32'b01111111111111100000000000000000;
			13'h1087: data = 32'b01111111111111111110000000000000;
			13'h1088: data = 32'b01111111111111111111100000000000;
			13'h1089: data = 32'b01111111111111111111110000000000;
			13'h108a: data = 32'b00111111111111111111111000000000;
			13'h108b: data = 32'b00000111111111111111111000000000;
			13'h108c: data = 32'b00000111111000001111111100000000;
			13'h108d: data = 32'b00000111111000000011111100000000;
			13'h108e: data = 32'b00000111111000000011111110000000;
			13'h108f: data = 32'b00000111111000000001111110000000;
			13'h1090: data = 32'b00000111111000000001111110000000;
			13'h1091: data = 32'b00000111111000000001111110000000;
			13'h1092: data = 32'b00000111111000000001111110000000;
			13'h1093: data = 32'b00000111111000000001111110000000;
			13'h1094: data = 32'b00000111111000000001111110000000;
			13'h1095: data = 32'b00000111111000000001111110000000;
			13'h1096: data = 32'b00000111111000000001111110000000;
			13'h1097: data = 32'b00000111111000000001111110000000;
			13'h1098: data = 32'b00000111111000000001111110000000;
			13'h1099: data = 32'b00000111111000000011111110000000;
			13'h109a: data = 32'b00000111111000000011111100000000;
			13'h109b: data = 32'b00000111111000001111111100000000;
			13'h109c: data = 32'b00000111111111111111111000000000;
			13'h109d: data = 32'b00000111111111111111110000000000;
			13'h109e: data = 32'b00000111111111111111100000000000;
			13'h109f: data = 32'b00000111111111111111111000000000;
			13'h10a0: data = 32'b00000111111111111111111100000000;
			13'h10a1: data = 32'b00000111111000111111111100000000;
			13'h10a2: data = 32'b00000111111000000111111110000000;
			13'h10a3: data = 32'b00000111111000000011111110000000;
			13'h10a4: data = 32'b00000111111000000001111111000000;
			13'h10a5: data = 32'b00000111111000000001111111000000;
			13'h10a6: data = 32'b00000111111000000000111111000000;
			13'h10a7: data = 32'b00000111111000000000111111100000;
			13'h10a8: data = 32'b00000111111000000000111111100000;
			13'h10a9: data = 32'b00000111111000000000111111100000;
			13'h10aa: data = 32'b00000111111000000000111111100000;
			13'h10ab: data = 32'b00000111111000000000111111100000;
			13'h10ac: data = 32'b00000111111000000000111111100000;
			13'h10ad: data = 32'b00000111111000000000111111100000;
			13'h10ae: data = 32'b00000111111000000000111111000000;
			13'h10af: data = 32'b00000111111000000000111111000000;
			13'h10b0: data = 32'b00000111111000000001111111000000;
			13'h10b1: data = 32'b00000111111000000001111111000000;
			13'h10b2: data = 32'b00000111111000000111111110000000;
			13'h10b3: data = 32'b00000111111100011111111110000000;
			13'h10b4: data = 32'b00001111111111111111111100000000;
			13'h10b5: data = 32'b01111111111111111111111000000000;
			13'h10b6: data = 32'b01111111111111111111110000000000;
			13'h10b7: data = 32'b01111111111111111111100000000000;
			13'h10b8: data = 32'b01111111111111111110000000000000;
			13'h10b9: data = 32'b00000000000000000000000000000000;
			13'h10ba: data = 32'b00000000000000000000000000000000;
			13'h10bb: data = 32'b00000000000000000000000000000000;
			13'h10bc: data = 32'b00000000000000000000000000000000;
			13'h10bd: data = 32'b00000000000000000000000000000000;
			13'h10be: data = 32'b00000000000000000000000000000000;
			13'h10bf: data = 32'b00000000000000000000000000000000;
//C x4
			13'h10c0: data = 32'b00000000000001111111111000000000;
			13'h10c1: data = 32'b00000000000011111111111100000000;
			13'h10c2: data = 32'b00000000001111111111111110000000;
			13'h10c3: data = 32'b00000000011111111111111111000000;
			13'h10c4: data = 32'b00000000111111111111111111100000;
			13'h10c5: data = 32'b00000000111111111111111111110000;
			13'h10c6: data = 32'b00000001111111111111111111110000;
			13'h10c7: data = 32'b00000011111111111111111111111000;
			13'h10c8: data = 32'b00000011111111111111111111111000;
			13'h10c9: data = 32'b00000111111111100000011111111100;
			13'h10ca: data = 32'b00000111111111000000001111111100;
			13'h10cb: data = 32'b00000111111110000000000111111110;
			13'h10cc: data = 32'b00001111111100000000000111111110;
			13'h10cd: data = 32'b00001111111100000000000011111110;
			13'h10ce: data = 32'b00001111111000000000000011111110;
			13'h10cf: data = 32'b00011111111000000000000001111111;
			13'h10d0: data = 32'b00011111110000000000000001111111;
			13'h10d1: data = 32'b00011111110000000000000001111111;
			13'h10d2: data = 32'b00011111110000000000000001111111;
			13'h10d3: data = 32'b00011111110000000000000001111111;
			13'h10d4: data = 32'b00011111100000000000000000111000;
			13'h10d5: data = 32'b00111111100000000000000000000000;
			13'h10d6: data = 32'b00111111100000000000000000000000;
			13'h10d7: data = 32'b00111111100000000000000000000000;
			13'h10d8: data = 32'b00111111100000000000000000000000;
			13'h10d9: data = 32'b00111111100000000000000000000000;
			13'h10da: data = 32'b00111111100000000000000000000000;
			13'h10db: data = 32'b00111111100000000000000000000000;
			13'h10dc: data = 32'b00111111100000000000000000000000;
			13'h10dd: data = 32'b00111111100000000000000000000000;
			13'h10de: data = 32'b00111111100000000000000000000000;
			13'h10df: data = 32'b00111111100000000000000000000000;
			13'h10e0: data = 32'b00111111100000000000000000000000;
			13'h10e1: data = 32'b00111111100000000000000000000000;
			13'h10e2: data = 32'b00111111100000000000000000000000;
			13'h10e3: data = 32'b00111111100000000000000000000000;
			13'h10e4: data = 32'b00111111100000000000000000000000;
			13'h10e5: data = 32'b00111111100000000000000000000000;
			13'h10e6: data = 32'b00111111100000000000000000000000;
			13'h10e7: data = 32'b00111111100000000000000000000000;
			13'h10e8: data = 32'b00111111100000000000000000111000;
			13'h10e9: data = 32'b00111111100000000000000000111111;
			13'h10ea: data = 32'b00111111100000000000000000111111;
			13'h10eb: data = 32'b00111111100000000000000000111111;
			13'h10ec: data = 32'b00011111110000000000000000111111;
			13'h10ed: data = 32'b00011111110000000000000001111111;
			13'h10ee: data = 32'b00011111110000000000000001111111;
			13'h10ef: data = 32'b00011111110000000000000001111111;
			13'h10f0: data = 32'b00011111111000000000000001111111;
			13'h10f1: data = 32'b00001111111000000000000011111110;
			13'h10f2: data = 32'b00001111111000000000000011111110;
			13'h10f3: data = 32'b00001111111100000000000111111110;
			13'h10f4: data = 32'b00000111111110000000000111111100;
			13'h10f5: data = 32'b00000111111111000000001111111100;
			13'h10f6: data = 32'b00000111111111100000011111111100;
			13'h10f7: data = 32'b00000011111111111111111111111000;
			13'h10f8: data = 32'b00000011111111111111111111111000;
			13'h10f9: data = 32'b00000001111111111111111111110000;
			13'h10fa: data = 32'b00000000111111111111111111110000;
			13'h10fb: data = 32'b00000000111111111111111111100000;
			13'h10fc: data = 32'b00000000011111111111111111000000;
			13'h10fd: data = 32'b00000000001111111111111110000000;
			13'h10fe: data = 32'b00000000000111111111111100000000;
			13'h10ff: data = 32'b00000000000001111111110000000000;
			  
// D x44
			13'h1100: data = 32'b00000000000000000000000000000000;
			13'h1101: data = 32'b00000000000000000000000000000000;
			13'h1102: data = 32'b00000000000000000000000000000000;
			13'h1103: data = 32'b00000000000000000000000000000000;
			13'h1104: data = 32'b00000000000000000000000000000000;
			13'h1105: data = 32'b00000111111111111110000000000000;
			13'h1106: data = 32'b00000111111111111111110000000000;
			13'h1107: data = 32'b00000111111111111111111000000000;
			13'h1108: data = 32'b00000111111111111111111100000000;
			13'h1109: data = 32'b00000111111111111111111110000000;
			13'h110a: data = 32'b00000111111111111111111110000000;
			13'h110b: data = 32'b00000111111111111111111111000000;
			13'h110c: data = 32'b00000111111111111111111111000000;
			13'h110d: data = 32'b00000111111111111111111111100000;
			13'h110e: data = 32'b00000111111111111111111111100000;
			13'h110f: data = 32'b00000111111111111111111111110000;
			13'h1110: data = 32'b00000111111100000001111111110000;
			13'h1111: data = 32'b00000111111100000000111111110000;
			13'h1112: data = 32'b00000111111100000000011111110000;
			13'h1113: data = 32'b00000111111100000000011111111000;
			13'h1114: data = 32'b00000111111100000000001111111000;
			13'h1115: data = 32'b00000111111100000000001111111000;
			13'h1116: data = 32'b00000111111100000000001111111000;
			13'h1117: data = 32'b00000111111100000000000111111000;
			13'h1118: data = 32'b00000111111100000000000111111000;
			13'h1119: data = 32'b00000111111100000000000111111000;
			13'h111a: data = 32'b00000111111100000000000111111100;
			13'h111b: data = 32'b00000111111100000000000111111100;
			13'h111c: data = 32'b00000111111100000000000111111100;
			13'h111d: data = 32'b00000111111100000000000111111100;
			13'h111e: data = 32'b00000111111100000000000111111100;
			13'h111f: data = 32'b00000111111100000000000111111100;
			13'h1120: data = 32'b00000111111100000000000111111100;
			13'h1121: data = 32'b00000111111100000000000111111100;
			13'h1122: data = 32'b00000111111100000000000111111100;
			13'h1123: data = 32'b00000111111100000000000111111100;
			13'h1124: data = 32'b00000111111100000000000111111100;
			13'h1125: data = 32'b00000111111100000000000111111100;
			13'h1126: data = 32'b00000111111100000000000111111100;
			13'h1127: data = 32'b00000111111100000000000111111100;
			13'h1128: data = 32'b00000111111100000000000111111100;
			13'h1129: data = 32'b00000111111100000000000111111100;
			13'h112a: data = 32'b00000111111100000000000111111000;
			13'h112b: data = 32'b00000111111100000000000111111000;
			13'h112c: data = 32'b00000111111100000000000111111000;
			13'h112d: data = 32'b00000111111100000000001111111000;
			13'h112e: data = 32'b00000111111100000000001111111000;
			13'h112f: data = 32'b00000111111100000000001111111000;
			13'h1130: data = 32'b00000111111100000000001111111000;
			13'h1131: data = 32'b00000111111100000000011111110000;
			13'h1132: data = 32'b00000111111100000000011111110000;
			13'h1133: data = 32'b00000111111100000000111111110000;
			13'h1134: data = 32'b00000111111111111111111111110000;
			13'h1135: data = 32'b00000111111111111111111111100000;
			13'h1136: data = 32'b00000111111111111111111111100000;
			13'h1137: data = 32'b00000111111111111111111111000000;
			13'h1138: data = 32'b00000111111111111111111111000000;
			13'h1139: data = 32'b00000111111111111111111110000000;
			13'h113a: data = 32'b00000111111111111111111110000000;
			13'h113b: data = 32'b00000111111111111111111100000000;
			13'h113c: data = 32'b00000111111111111111111000000000;
			13'h113d: data = 32'b00000111111111111111100000000000;
			13'h113e: data = 32'b00000111111111111100000000000000;
			13'h113f: data = 32'b00000000000000000000000000000000;

//E  x45
			13'h1140: data = 32'b00000001000000000000000000110000;
			13'h1141: data = 32'b00000011111111111111111111110000;
			13'h1142: data = 32'b00000011111111111111111111110000;
			13'h1143: data = 32'b00000011111111111111111111110000;
			13'h1144: data = 32'b00000011111111111111111111110000;
			13'h1145: data = 32'b00000011111111111111111111110000;
			13'h1146: data = 32'b00000011111111111111111111110000;
			13'h1147: data = 32'b00000011111111111111111111110000;
			13'h1148: data = 32'b00000011111111111111111111110000;
			13'h1149: data = 32'b00000011111111111111111111110000;
			13'h114a: data = 32'b00000011111111111111111111110000;
			13'h114b: data = 32'b00000011111111111111111111110000;
			13'h114c: data = 32'b00000011111111111111111111110000;
			13'h114d: data = 32'b00000011111111111111111111110000;
			13'h114e: data = 32'b00000011111111110000000000000000;
			13'h114f: data = 32'b00000011111111110000000000000000;
			13'h1150: data = 32'b00000011111111110000000000000000;
			13'h1151: data = 32'b00000011111111110000000000000000;
			13'h1152: data = 32'b00000011111111110000000000000000;
			13'h1153: data = 32'b00000011111111110000000000000000;
			13'h1154: data = 32'b00000011111111110000000000000000;
			13'h1155: data = 32'b00000011111111110000000000000000;
			13'h1156: data = 32'b00000011111111110000000000000000;
			13'h1157: data = 32'b00000011111111110000000000000000;
			13'h1158: data = 32'b00000011111111111111111111000000;
			13'h1159: data = 32'b00000011111111111111111111000000;
			13'h115a: data = 32'b00000011111111111111111111000000;
			13'h115b: data = 32'b00000011111111111111111111000000;
			13'h115c: data = 32'b00000011111111111111111111000000;
			13'h115d: data = 32'b00000011111111111111111111000000;
			13'h115e: data = 32'b00000011111111111111111111000000;
			13'h115f: data = 32'b00000011111111111111111111000000;
			13'h1160: data = 32'b00000011111111111111111111000000;
			13'h1161: data = 32'b00000011111111111111111111000000;
			13'h1162: data = 32'b00000011111111111111111111000000;
			13'h1163: data = 32'b00000011111111111111111111000000;
			13'h1164: data = 32'b00000011111111110000000000000000;
			13'h1165: data = 32'b00000011111111110000000000000000;
			13'h1166: data = 32'b00000011111111110000000000000000;
			13'h1167: data = 32'b00000011111111110000000000000000;
			13'h1168: data = 32'b00000011111111110000000000000000;
			13'h1169: data = 32'b00000011111111110000000000000000;
			13'h116a: data = 32'b00000011111111110000000000000000;
			13'h116b: data = 32'b00000011111111110000000000000000;
			13'h116c: data = 32'b00000011111111110000000000000000;
			13'h116d: data = 32'b00000011111111110000000000000000;
			13'h116e: data = 32'b00000011111111110000000000000000;
			13'h116f: data = 32'b00000011111111110000000000000000;
			13'h1170: data = 32'b00000011111111111111111111110000;
			13'h1171: data = 32'b00000011111111111111111111110000;
			13'h1172: data = 32'b00000011111111111111111111110000;
			13'h1173: data = 32'b00000011111111111111111111110000;
			13'h1174: data = 32'b00000011111111111111111111110000;
			13'h1175: data = 32'b00000011111111111111111111110000;
			13'h1176: data = 32'b00000011111111111111111111110000;
			13'h1177: data = 32'b00000011111111111111111111110000;
			13'h1178: data = 32'b00000011111111111111111111110000;
			13'h1179: data = 32'b00000011111111111111111111110000;
			13'h117a: data = 32'b00000011111111111111111111110000;
			13'h117b: data = 32'b00000011111111111111111111110000;
			13'h117c: data = 32'b00000011111111111111111111110000;
			13'h117d: data = 32'b00000000000000000000000000000000;
			13'h117e: data = 32'b00000000000000000000000000000000;
			13'h117f: data = 32'b00000000000000000000000000000000;

// F x46
			13'h1180: data = 32'b00000000000000000000000000000000;
			13'h1181: data = 32'b00000000000000000000000000000000;
			13'h1182: data = 32'b00000000000000000000000000000000;
			13'h1183: data = 32'b00000000000000000000000000000000;
			13'h1184: data = 32'b01111111111111111111111111110000;
			13'h1185: data = 32'b01111111111111111111111111111000;
			13'h1186: data = 32'b01111111111111111111111111111000;
			13'h1187: data = 32'b01111111111111111111111111111000;
			13'h1188: data = 32'b00111111111111111111111111111000;
			13'h1189: data = 32'b00001111111111111111111111111000;
			13'h118a: data = 32'b00000111111100000000000111111000;
			13'h118b: data = 32'b00000111111100000000000011111000;
			13'h118c: data = 32'b00000111111100000000000001111000;
			13'h118d: data = 32'b00000111111100000000000001111000;
			13'h118e: data = 32'b00000111111100000000000001111000;
			13'h118f: data = 32'b00000111111100000000000001111000;
			13'h1190: data = 32'b00000111111100000000000001111000;
			13'h1191: data = 32'b00000111111100000000000001111000;
			13'h1192: data = 32'b00000111111100000000000000111000;
			13'h1193: data = 32'b00000111111100000000000000000000;
			13'h1194: data = 32'b00000111111100000000001110000000;
			13'h1195: data = 32'b00000111111100000000001110000000;
			13'h1196: data = 32'b00000111111100000000001110000000;
			13'h1197: data = 32'b00000111111100000000001110000000;
			13'h1198: data = 32'b00000111111100000000001110000000;
			13'h1199: data = 32'b00000111111100000000001110000000;
			13'h119a: data = 32'b00000111111100000000011110000000;
			13'h119b: data = 32'b00000111111100000000111110000000;
			13'h119c: data = 32'b00000111111111111111111110000000;
			13'h119d: data = 32'b00000111111111111111111110000000;
			13'h119e: data = 32'b00000111111111111111111110000000;
			13'h119f: data = 32'b00000111111111111111111110000000;
			13'h11a0: data = 32'b00000111111111111111111110000000;
			13'h11a1: data = 32'b00000111111111111111111110000000;
			13'h11a2: data = 32'b00000111111100000000111110000000;
			13'h11a3: data = 32'b00000111111100000000011110000000;
			13'h11a4: data = 32'b00000111111100000000001110000000;
			13'h11a5: data = 32'b00000111111100000000001110000000;
			13'h11a6: data = 32'b00000111111100000000001110000000;
			13'h11a7: data = 32'b00000111111100000000001110000000;
			13'h11a8: data = 32'b00000111111100000000001110000000;
			13'h11a9: data = 32'b00000111111100000000001110000000;
			13'h11aa: data = 32'b00000111111100000000000000000000;
			13'h11ab: data = 32'b00000111111100000000000000000000;
			13'h11ac: data = 32'b00000111111100000000000000000000;
			13'h11ad: data = 32'b00000111111100000000000000000000;
			13'h11ae: data = 32'b00000111111100000000000000000000;
			13'h11af: data = 32'b00000111111100000000000000000000;
			13'h11b0: data = 32'b00000111111100000000000000000000;
			13'h11b1: data = 32'b00000111111100000000000000000000;
			13'h11b2: data = 32'b00000111111100000000000000000000;
			13'h11b3: data = 32'b00000111111100000000000000000000;
			13'h11b4: data = 32'b00000111111100000000000000000000;
			13'h11b5: data = 32'b00000111111100000000000000000000;
			13'h11b6: data = 32'b00000111111100000000000000000000;
			13'h11b7: data = 32'b00001111111110000000000000000000;
			13'h11b8: data = 32'b01111111111111110000000000000000;
			13'h11b9: data = 32'b01111111111111110000000000000000;
			13'h11ba: data = 32'b01111111111111110000000000000000;
			13'h11bb: data = 32'b01111111111111110000000000000000;
			13'h11bc: data = 32'b01111111111111110000000000000000;
			13'h11bd: data = 32'b00000000000000000000000000000000;
			13'h11be: data = 32'b00000000000000000000000000000000;
			13'h11bf: data = 32'b00000000000000000000000000000000;

//G x47
			13'h11c0: data = 32'b00000000000000000000000000000000;
			13'h11c1: data = 32'b00000000000000000000000000000000;
			13'h11c2: data = 32'b00000000000000000000000000000000;
			13'h11c3: data = 32'b00000000000000000000000000000000;
			13'h11c4: data = 32'b00000000000000000000000000000000;
			13'h11c5: data = 32'b00000000000000000000000000000000;
			13'h11c6: data = 32'b00000000000000000000000000000000;
			13'h11c7: data = 32'b00000000000000111111000000000000;
			13'h11c8: data = 32'b00000000000001111111110000000000;
			13'h11c9: data = 32'b00000000000011111111111000000000;
			13'h11ca: data = 32'b00000000000111111111111000000000;
			13'h11cb: data = 32'b00000000001111111111111100000000;
			13'h11cc: data = 32'b00000000001111111111111100000000;
			13'h11cd: data = 32'b00000000011111110011111110000000;
			13'h11ce: data = 32'b00000000011111000000111110000000;
			13'h11cf: data = 32'b00000000111110000000011110000000;
			13'h11d0: data = 32'b00000000111110000000011111000000;
			13'h11d1: data = 32'b00000000111100000000001111000000;
			13'h11d2: data = 32'b00000001111100000000001111000000;
			13'h11d3: data = 32'b00000001111000000000001111000000;
			13'h11d4: data = 32'b00000001111000000000001111000000;
			13'h11d5: data = 32'b00000001111000000000000111000000;
			13'h11d6: data = 32'b00000001111000000000000111000000;
			13'h11d7: data = 32'b00000001110000000000000110000000;
			13'h11d8: data = 32'b00000011110000000000000000000000;
			13'h11d9: data = 32'b00000011110000000000000000000000;
			13'h11da: data = 32'b00000011110000000000000000000000;
			13'h11db: data = 32'b00000011110000000000000000000000;
			13'h11dc: data = 32'b00000011110000000000000000000000;
			13'h11dd: data = 32'b00000011110000000000000000000000;
			13'h11de: data = 32'b00000011110000000000000000000000;
			13'h11df: data = 32'b00000011110000000000000000000000;
			13'h11e0: data = 32'b00000011110000000000000000000000;
			13'h11e1: data = 32'b00000011110000000111111111100000;
			13'h11e2: data = 32'b00000011110000000111111111100000;
			13'h11e3: data = 32'b00000011110000000111111111100000;
			13'h11e4: data = 32'b00000011110000000111111111100000;
			13'h11e5: data = 32'b00000011110000000111111111100000;
			13'h11e6: data = 32'b00000011110000000111111111100000;
			13'h11e7: data = 32'b00000011110000000111111111100000;
			13'h11e8: data = 32'b00000011110000000000000111100000;
			13'h11e9: data = 32'b00000011110000000000000111100000;
			13'h11ea: data = 32'b00000011110000000000000111100000;
			13'h11eb: data = 32'b00000001110000000000000111100000;
			13'h11ec: data = 32'b00000001111000000000000111100000;
			13'h11ed: data = 32'b00000001111000000000000111100000;
			13'h11ee: data = 32'b00000001111000000000000111100000;
			13'h11ef: data = 32'b00000001111000000000000111100000;
			13'h11f0: data = 32'b00000001111100000000000111100000;
			13'h11f1: data = 32'b00000000111100000000000111100000;
			13'h11f2: data = 32'b00000000111110000000001111100000;
			13'h11f3: data = 32'b00000000111111000000011111100000;
			13'h11f4: data = 32'b00000000011111100000111111100000;
			13'h11f5: data = 32'b00000000011111111111111111000000;
			13'h11f6: data = 32'b00000000001111111111111110000000;
			13'h11f7: data = 32'b00000000001111111111111110000000;
			13'h11f8: data = 32'b00000000000111111111111100000000;
			13'h11f9: data = 32'b00000000000011111111111000000000;
			13'h11fa: data = 32'b00000000000001111111110000000000;
			13'h11fb: data = 32'b00000000000000111111100000000000;
			13'h11fc: data = 32'b00000000000000000000000000000000;
			13'h11fd: data = 32'b00000000000000000000000000000000;
			13'h11fe: data = 32'b00000000000000000000000000000000;
			13'h11ff: data = 32'b00000000000000000000000000000000;


//H x48
			13'h1200: data = 32'b00000000000000000000000000000000;
			13'h1201: data = 32'b00111111100000000000011111110000;
			13'h1202: data = 32'b00111111100000000000011111110000;
			13'h1203: data = 32'b00111111100000000000011111110000;
			13'h1204: data = 32'b00111111100000000000011111110000;
			13'h1205: data = 32'b00111111100000000000011111110000;
			13'h1206: data = 32'b00111111100000000000011111110000;
			13'h1207: data = 32'b00111111100000000000011111110000;
			13'h1208: data = 32'b00111111100000000000011111110000;
			13'h1209: data = 32'b00111111100000000000011111110000;
			13'h120a: data = 32'b00111111100000000000011111110000;
			13'h120b: data = 32'b00111111100000000000011111110000;
			13'h120c: data = 32'b00111111100000000000011111110000;
			13'h120d: data = 32'b00111111100000000000011111110000;
			13'h120e: data = 32'b00111111100000000000011111110000;
			13'h120f: data = 32'b00111111100000000000011111110000;
			13'h1210: data = 32'b00111111100000000000011111110000;
			13'h1211: data = 32'b00111111100000000000011111110000;
			13'h1212: data = 32'b00111111100000000000011111110000;
			13'h1213: data = 32'b00111111100000000000011111110000;
			13'h1214: data = 32'b00111111100000000000011111110000;
			13'h1215: data = 32'b00111111100000000000011111110000;
			13'h1216: data = 32'b00111111100000000000011111110000;
			13'h1217: data = 32'b00111111100000000000011111110000;
			13'h1218: data = 32'b00111111100000000000011111110000;
			13'h1219: data = 32'b00111111111111111111111111110000;
			13'h121a: data = 32'b00111111111111111111111111110000;
			13'h121b: data = 32'b00111111111111111111111111110000;
			13'h121c: data = 32'b00111111111111111111111111110000;
			13'h121d: data = 32'b00111111111111111111111111110000;
			13'h121e: data = 32'b00111111111111111111111111110000;
			13'h121f: data = 32'b00111111111111111111111111110000;
			13'h1220: data = 32'b00111111111111111111111111110000;
			13'h1221: data = 32'b00111111111111111111111111110000;
			13'h1222: data = 32'b00111111111111111111111111110000;
			13'h1223: data = 32'b00111111111111111111111111110000;
			13'h1224: data = 32'b00111111100000000000011111110000;
			13'h1225: data = 32'b00111111100000000000011111110000;
			13'h1226: data = 32'b00111111100000000000011111110000;
			13'h1227: data = 32'b00111111100000000000011111110000;
			13'h1228: data = 32'b00111111100000000000011111110000;
			13'h1229: data = 32'b00111111100000000000011111110000;
			13'h122a: data = 32'b00111111100000000000011111110000;
			13'h122b: data = 32'b00111111100000000000011111110000;
			13'h122c: data = 32'b00111111100000000000011111110000;
			13'h122d: data = 32'b00111111100000000000011111110000;
			13'h122e: data = 32'b00111111100000000000011111110000;
			13'h122f: data = 32'b00111111100000000000011111110000;
			13'h1230: data = 32'b00111111100000000000011111110000;
			13'h1231: data = 32'b00111111100000000000011111110000;
			13'h1232: data = 32'b00111111100000000000011111110000;
			13'h1233: data = 32'b00111111100000000000011111110000;
			13'h1234: data = 32'b00111111100000000000011111110000;
			13'h1235: data = 32'b00111111100000000000011111110000;
			13'h1236: data = 32'b00111111100000000000011111110000;
			13'h1237: data = 32'b00111111100000000000011111110000;
			13'h1238: data = 32'b00111111100000000000011111110000;
			13'h1239: data = 32'b00111111100000000000011111110000;
			13'h123a: data = 32'b00111111100000000000011111110000;
			13'h123b: data = 32'b00111111100000000000011111110000;
			13'h123c: data = 32'b00111111100000000000011111110000;
			13'h123d: data = 32'b00111111100000000000011111110000;
			13'h123e: data = 32'b00000000000000000000000000000000;
			13'h123f: data = 32'b00000000000000000000000000000000;

//I x49
			13'h1240: data = 32'b00000000000000000000000000000000;
			13'h1241: data = 32'b00001111111111111111111100000000;
			13'h1242: data = 32'b00001111111111111111111100000000;
			13'h1243: data = 32'b00001111111111111111111100000000;
			13'h1244: data = 32'b00001111111111111111111100000000;
			13'h1245: data = 32'b00001111111111111111111100000000;
			13'h1246: data = 32'b00001111111111111111111100000000;
			13'h1247: data = 32'b00001111111111111111111100000000;
			13'h1248: data = 32'b00001111111111111111111100000000;
			13'h1249: data = 32'b00001111111111111111111100000000;
			13'h124a: data = 32'b00000111101111111111111000000000;
			13'h124b: data = 32'b00000000001111111100000000000000;
			13'h124c: data = 32'b00000000001111111100000000000000;
			13'h124d: data = 32'b00000000001111111100000000000000;
			13'h124e: data = 32'b00000000001111111100000000000000;
			13'h124f: data = 32'b00000000001111111100000000000000;
			13'h1250: data = 32'b00000000001111111100000000000000;
			13'h1251: data = 32'b00000000001111111100000000000000;
			13'h1252: data = 32'b00000000001111111100000000000000;
			13'h1253: data = 32'b00000000001111111100000000000000;
			13'h1254: data = 32'b00000000001111111100000000000000;
			13'h1255: data = 32'b00000000001111111100000000000000;
			13'h1256: data = 32'b00000000001111111100000000000000;
			13'h1257: data = 32'b00000000001111111100000000000000;
			13'h1258: data = 32'b00000000001111111100000000000000;
			13'h1259: data = 32'b00000000001111111100000000000000;
			13'h125a: data = 32'b00000000001111111100000000000000;
			13'h125b: data = 32'b00000000001111111100000000000000;
			13'h125c: data = 32'b00000000001111111100000000000000;
			13'h125d: data = 32'b00000000001111111100000000000000;
			13'h125e: data = 32'b00000000001111111100000000000000;
			13'h125f: data = 32'b00000000001111111100000000000000;
			13'h1260: data = 32'b00000000001111111100000000000000;
			13'h1261: data = 32'b00000000001111111100000000000000;
			13'h1262: data = 32'b00000000001111111100000000000000;
			13'h1263: data = 32'b00000000001111111100000000000000;
			13'h1264: data = 32'b00000000001111111100000000000000;
			13'h1265: data = 32'b00000000001111111100000000000000;
			13'h1266: data = 32'b00000000001111111100000000000000;
			13'h1267: data = 32'b00000000001111111100000000000000;
			13'h1268: data = 32'b00000000001111111100000000000000;
			13'h1269: data = 32'b00000000001111111100000000000000;
			13'h126a: data = 32'b00000000001111111100000000000000;
			13'h126b: data = 32'b00000000001111111100000000000000;
			13'h126c: data = 32'b00000000001111111100000000000000;
			13'h126d: data = 32'b00000000001111111100000000000000;
			13'h126e: data = 32'b00000000001111111100000000000000;
			13'h126f: data = 32'b00000000001111111100000000000000;
			13'h1270: data = 32'b00000000001111111100000000000000;
			13'h1271: data = 32'b00000000001111111100000000000000;
			13'h1272: data = 32'b00000000001111111100000000000000;
			13'h1273: data = 32'b00000000001111111100000000000000;
			13'h1274: data = 32'b00000000001111111100000000000000;
			13'h1275: data = 32'b00000111111111111111111100000000;
			13'h1276: data = 32'b00001111111111111111111100000000;
			13'h1277: data = 32'b00001111111111111111111100000000;
			13'h1278: data = 32'b00001111111111111111111100000000;
			13'h1279: data = 32'b00001111111111111111111100000000;
			13'h127a: data = 32'b00001111111111111111111100000000;
			13'h127b: data = 32'b00001111111111111111111100000000;
			13'h127c: data = 32'b00001111111111111111111100000000;
			13'h127d: data = 32'b00001111111111111111111100000000;
			13'h127e: data = 32'b00001111111111111111111100000000;
			13'h127f: data = 32'b00000000000000000000000000000000;


//J x4a
			13'h1280: data = 32'b00000000000000000000000000000000;
			13'h1281: data = 32'b00000000000000000000011111111100;
			13'h1282: data = 32'b00000000000000000000011111111100;
			13'h1283: data = 32'b00000000000000000000011111111100;
			13'h1284: data = 32'b00000000000000000000011111111100;
			13'h1285: data = 32'b00000000000000000000011111111100;
			13'h1286: data = 32'b00000000000000000000011111111100;
			13'h1287: data = 32'b00000000000000000000011111111100;
			13'h1288: data = 32'b00000000000000000000011111111100;
			13'h1289: data = 32'b00000000000000000000011111111100;
			13'h128a: data = 32'b00000000000000000000011111111100;
			13'h128b: data = 32'b00000000000000000000011111111100;
			13'h128c: data = 32'b00000000000000000000011111111100;
			13'h128d: data = 32'b00000000000000000000011111111100;
			13'h128e: data = 32'b00000000000000000000011111111100;
			13'h128f: data = 32'b00000000000000000000011111111100;
			13'h1290: data = 32'b00000000000000000000011111111100;
			13'h1291: data = 32'b00000000000000000000011111111100;
			13'h1292: data = 32'b00000000000000000000011111111100;
			13'h1293: data = 32'b00000000000000000000011111111100;
			13'h1294: data = 32'b00000000000000000000011111111100;
			13'h1295: data = 32'b00000000000000000000011111111100;
			13'h1296: data = 32'b00000000000000000000011111111100;
			13'h1297: data = 32'b00000000000000000000011111111100;
			13'h1298: data = 32'b00000000000000000000011111111100;
			13'h1299: data = 32'b00000000000000000000011111111100;
			13'h129a: data = 32'b00000000000000000000011111111100;
			13'h129b: data = 32'b00000000000000000000011111111100;
			13'h129c: data = 32'b00000000000000000000011111111100;
			13'h129d: data = 32'b00000000000000000000011111111100;
			13'h129e: data = 32'b00000000000000000000011111111100;
			13'h129f: data = 32'b00000000000000000000011111111100;
			13'h12a0: data = 32'b00000000000000000000011111111100;
			13'h12a1: data = 32'b00000000000000000000011111111100;
			13'h12a2: data = 32'b00000000000000000000011111111100;
			13'h12a3: data = 32'b00000000000000000000011111111100;
			13'h12a4: data = 32'b00000000000000000000011111111100;
			13'h12a5: data = 32'b00000000000000000000011111111100;
			13'h12a6: data = 32'b00000000000000000000011111111100;
			13'h12a7: data = 32'b00000000000000000000011111111100;
			13'h12a8: data = 32'b00000000000000000000011111111100;
			13'h12a9: data = 32'b00000000111000000000011111111100;
			13'h12aa: data = 32'b00111111111000000000011111111100;
			13'h12ab: data = 32'b00111111111000000000011111111100;
			13'h12ac: data = 32'b00111111111000000000111111111100;
			13'h12ad: data = 32'b00111111111000000000111111111100;
			13'h12ae: data = 32'b00111111111000000000111111111100;
			13'h12af: data = 32'b00111111111100000000111111111100;
			13'h12b0: data = 32'b00011111111100000000111111111000;
			13'h12b1: data = 32'b00011111111100000000111111111000;
			13'h12b2: data = 32'b00011111111110000001111111111000;
			13'h12b3: data = 32'b00011111111111100111111111111000;
			13'h12b4: data = 32'b00011111111111111111111111111000;
			13'h12b5: data = 32'b00001111111111111111111111110000;
			13'h12b6: data = 32'b00001111111111111111111111110000;
			13'h12b7: data = 32'b00001111111111111111111111100000;
			13'h12b8: data = 32'b00000111111111111111111111100000;
			13'h12b9: data = 32'b00000011111111111111111111000000;
			13'h12ba: data = 32'b00000011111111111111111110000000;
			13'h12bb: data = 32'b00000001111111111111111100000000;
			13'h12bc: data = 32'b00000000111111111111111000000000;
			13'h12bd: data = 32'b00000000001111111111110000000000;
			13'h12be: data = 32'b00000000000011111110000000000000;
			13'h12bf: data = 32'b00000000000000000000000000000000;

//K x4b
			13'h12c0: data = 32'b00000000000000000000000000000000;
			13'h12c1: data = 32'b01111111000000000000111111110000;
			13'h12c2: data = 32'b01111111000000000001111111110000;
			13'h12c3: data = 32'b01111111000000000001111111100000;
			13'h12c4: data = 32'b01111111000000000011111111100000;
			13'h12c5: data = 32'b01111111000000000011111111000000;
			13'h12c6: data = 32'b01111111000000000111111111000000;
			13'h12c7: data = 32'b01111111000000000111111110000000;
			13'h12c8: data = 32'b01111111000000001111111110000000;
			13'h12c9: data = 32'b01111111000000001111111100000000;
			13'h12ca: data = 32'b01111111000000011111111100000000;
			13'h12cb: data = 32'b01111111000000011111111000000000;
			13'h12cc: data = 32'b01111111000000111111111000000000;
			13'h12cd: data = 32'b01111111000000111111110000000000;
			13'h12ce: data = 32'b01111111000001111111110000000000;
			13'h12cf: data = 32'b01111111000001111111100000000000;
			13'h12d0: data = 32'b01111111000011111111100000000000;
			13'h12d1: data = 32'b01111111000011111111000000000000;
			13'h12d2: data = 32'b01111111000111111111000000000000;
			13'h12d3: data = 32'b01111111000111111110000000000000;
			13'h12d4: data = 32'b01111111001111111110000000000000;
			13'h12d5: data = 32'b01111111001111111100000000000000;
			13'h12d6: data = 32'b01111111011111111100000000000000;
			13'h12d7: data = 32'b01111111011111111000000000000000;
			13'h12d8: data = 32'b01111111111111111000000000000000;
			13'h12d9: data = 32'b01111111111111111000000000000000;
			13'h12da: data = 32'b01111111111111111000000000000000;
			13'h12db: data = 32'b01111111111111111000000000000000;
			13'h12dc: data = 32'b01111111111111111100000000000000;
			13'h12dd: data = 32'b01111111111111111100000000000000;
			13'h12de: data = 32'b01111111111111111110000000000000;
			13'h12df: data = 32'b01111111111111111110000000000000;
			13'h12e0: data = 32'b01111111111111111110000000000000;
			13'h12e1: data = 32'b01111111111111111111000000000000;
			13'h12e2: data = 32'b01111111111111111111000000000000;
			13'h12e3: data = 32'b01111111111001111111000000000000;
			13'h12e4: data = 32'b01111111111001111111100000000000;
			13'h12e5: data = 32'b01111111110001111111100000000000;
			13'h12e6: data = 32'b01111111110000111111100000000000;
			13'h12e7: data = 32'b01111111100000111111110000000000;
			13'h12e8: data = 32'b01111111100000111111110000000000;
			13'h12e9: data = 32'b01111111000000011111110000000000;
			13'h12ea: data = 32'b01111111000000011111111000000000;
			13'h12eb: data = 32'b01111111000000011111111000000000;
			13'h12ec: data = 32'b01111111000000001111111000000000;
			13'h12ed: data = 32'b01111111000000001111111100000000;
			13'h12ee: data = 32'b01111111000000001111111100000000;
			13'h12ef: data = 32'b01111111000000000111111100000000;
			13'h12f0: data = 32'b01111111000000000111111110000000;
			13'h12f1: data = 32'b01111111000000000111111110000000;
			13'h12f2: data = 32'b01111111000000000011111110000000;
			13'h12f3: data = 32'b01111111000000000011111111000000;
			13'h12f4: data = 32'b01111111000000000011111111000000;
			13'h12f5: data = 32'b01111111000000000001111111100000;
			13'h12f6: data = 32'b01111111000000000001111111100000;
			13'h12f7: data = 32'b01111111000000000001111111100000;
			13'h12f8: data = 32'b01111111000000000000111111110000;
			13'h12f9: data = 32'b01111111000000000000111111110000;
			13'h12fa: data = 32'b01111111000000000000111111110000;
			13'h12fb: data = 32'b01111111000000000000011111111000;
			13'h12fc: data = 32'b01111111000000000000011111111000;
			13'h12fd: data = 32'b01111111000000000000011111111000;
			13'h12fe: data = 32'b00000000000000000000000000000000;
			13'h12ff: data = 32'b00000000000000000000000000000000;

//L x4c
			13'h1300: data = 32'b00000000000000000000000000000000;
			13'h1301: data = 32'b00000000000000000000000000000000;
			13'h1302: data = 32'b01111111111111111110000000000000;
			13'h1303: data = 32'b01111111111111111110000000000000;
			13'h1304: data = 32'b01111111111111111110000000000000;
			13'h1305: data = 32'b01111111111111111110000000000000;
			13'h1306: data = 32'b01111111111111111110000000000000;
			13'h1307: data = 32'b01111111111111111110000000000000;
			13'h1308: data = 32'b01111111111111111110000000000000;
			13'h1309: data = 32'b01111111111111111110000000000000;
			13'h130a: data = 32'b01111111111111111110000000000000;
			13'h130b: data = 32'b01111111111111111110000000000000;
			13'h130c: data = 32'b01111111111111111110000000000000;
			13'h130d: data = 32'b01111111111111111110000000000000;
			13'h130e: data = 32'b01111111111111111110000000000000;
			13'h130f: data = 32'b00000011111111000000000000000000;
			13'h1310: data = 32'b00000011111111000000000000000000;
			13'h1311: data = 32'b00000011111111000000000000000000;
			13'h1312: data = 32'b00000011111111000000000000000000;
			13'h1313: data = 32'b00000011111111000000000000000000;
			13'h1314: data = 32'b00000011111111000000000000000000;
			13'h1315: data = 32'b00000011111111000000000000000000;
			13'h1316: data = 32'b00000011111111000000000000000000;
			13'h1317: data = 32'b00000011111111000000000000000000;
			13'h1318: data = 32'b00000011111111000000000000000000;
			13'h1319: data = 32'b00000011111111000000000000000000;
			13'h131a: data = 32'b00000011111111000000000000000000;
			13'h131b: data = 32'b00000011111111000000000000000000;
			13'h131c: data = 32'b00000011111111000000000000000000;
			13'h131d: data = 32'b00000011111111000000000000000000;
			13'h131e: data = 32'b00000011111111000000000000000000;
			13'h131f: data = 32'b00000011111111000000000000000000;
			13'h1320: data = 32'b00000011111111000000000000000000;
			13'h1321: data = 32'b00000011111111000000000000000000;
			13'h1322: data = 32'b00000011111111000000000000000000;
			13'h1323: data = 32'b00000011111111000000000000000000;
			13'h1324: data = 32'b00000011111111000000000000000000;
			13'h1325: data = 32'b00000011111111000000000000000000;
			13'h1326: data = 32'b00000011111111000000000000000000;
			13'h1327: data = 32'b00000011111111000000000001000010;
			13'h1328: data = 32'b00000011111111000000000011111110;
			13'h1329: data = 32'b00000011111111000000000011111110;
			13'h132a: data = 32'b00000011111111000000000011111110;
			13'h132b: data = 32'b00000011111111000000000011111110;
			13'h132c: data = 32'b00000011111111000000000011111110;
			13'h132d: data = 32'b00000011111111000000000011111110;
			13'h132e: data = 32'b00000011111111000000000011111110;
			13'h132f: data = 32'b00000011111111000000000011111110;
			13'h1330: data = 32'b00000011111111000000000011111110;
			13'h1331: data = 32'b01111111111111111111111111111110;
			13'h1332: data = 32'b01111111111111111111111111111110;
			13'h1333: data = 32'b01111111111111111111111111111110;
			13'h1334: data = 32'b01111111111111111111111111111110;
			13'h1335: data = 32'b01111111111111111111111111111110;
			13'h1336: data = 32'b01111111111111111111111111111110;
			13'h1337: data = 32'b01111111111111111111111111111110;
			13'h1338: data = 32'b01111111111111111111111111111110;
			13'h1339: data = 32'b01111111111111111111111111111110;
			13'h133a: data = 32'b01111111111111111111111111111110;
			13'h133b: data = 32'b01111111111111111111111111111110;
			13'h133c: data = 32'b01111111111111111111111111111110;
			13'h133d: data = 32'b01111111111111111111111111111110;
			13'h133e: data = 32'b01111111111111111111111111111110;
			13'h133f: data = 32'b00000000000000000000000000000000;


//M x4d
			13'h1340: data = 32'b10000000000000000000000000000000;
			13'h1341: data = 32'b11111111100000000000000011111111;
			13'h1342: data = 32'b11111111100000000000000111111111;
			13'h1343: data = 32'b11111111100000000000000111111111;
			13'h1344: data = 32'b11111111100000000000000111111111;
			13'h1345: data = 32'b11111111100000000000000111111111;
			13'h1346: data = 32'b10111111110000000000000111111100;
			13'h1347: data = 32'b10011111110000000000001111111000;
			13'h1348: data = 32'b10011111110000000000001111111000;
			13'h1349: data = 32'b10011111110000000000001111111000;
			13'h134a: data = 32'b10011111110000000000001111111000;
			13'h134b: data = 32'b10011111110000000000001111111000;
			13'h134c: data = 32'b10011111111000000000001111111000;
			13'h134d: data = 32'b10011111111000000000011111111000;
			13'h134e: data = 32'b10011111111000000000011111111000;
			13'h134f: data = 32'b10011111111000000000011111111000;
			13'h1350: data = 32'b10011111111000000000011111111000;
			13'h1351: data = 32'b10011111111100000000011111111000;
			13'h1352: data = 32'b10011111111100000000111111111000;
			13'h1353: data = 32'b10011111111100000000111111111000;
			13'h1354: data = 32'b10011111111100000000111111111000;
			13'h1355: data = 32'b10011111111100000000111011111000;
			13'h1356: data = 32'b10011111111110000000111011111000;
			13'h1357: data = 32'b10011111111110000000111011111000;
			13'h1358: data = 32'b10011111111110000001111011111000;
			13'h1359: data = 32'b10011111111110000001111011111000;
			13'h135a: data = 32'b10011111111110000001111011111000;
			13'h135b: data = 32'b10011110111110000001110011111000;
			13'h135c: data = 32'b10011110111111000001110011111000;
			13'h135d: data = 32'b10011110111111000011110011111000;
			13'h135e: data = 32'b10011110111111000011110011111000;
			13'h135f: data = 32'b10011110111111000011110011111000;
			13'h1360: data = 32'b10011110111111000011110011111000;
			13'h1361: data = 32'b10011110011111100011100011111000;
			13'h1362: data = 32'b10011110011111100011100011111000;
			13'h1363: data = 32'b10011110011111100111100011111000;
			13'h1364: data = 32'b10011110011111100111100011111000;
			13'h1365: data = 32'b10011110011111100111100011111000;
			13'h1366: data = 32'b10011110001111100111000011111000;
			13'h1367: data = 32'b10011110001111110111000011111000;
			13'h1368: data = 32'b10011110001111111111000011111000;
			13'h1369: data = 32'b10011110001111111111000011111000;
			13'h136a: data = 32'b10011110001111111111000011111000;
			13'h136b: data = 32'b10011110000111111111000011111000;
			13'h136c: data = 32'b10011110000111111110000011111000;
			13'h136d: data = 32'b10011110000111111110000011111000;
			13'h136e: data = 32'b10011110000111111110000011111000;
			13'h136f: data = 32'b10011110000111111110000011111000;
			13'h1370: data = 32'b10011110000111111110000011111000;
			13'h1371: data = 32'b10011110000011111100000011111000;
			13'h1372: data = 32'b10011110000011111100000011111000;
			13'h1373: data = 32'b10011110000011111100000011111000;
			13'h1374: data = 32'b10011110000011111100000011111000;
			13'h1375: data = 32'b10011110000011111100000011111000;
			13'h1376: data = 32'b10011110000001111100000011111000;
			13'h1377: data = 32'b10011110000001111000000011111000;
			13'h1378: data = 32'b10011110000001111000000111111000;
			13'h1379: data = 32'b10111111000001111000000111111100;
			13'h137a: data = 32'b11111111110001111000011111111111;
			13'h137b: data = 32'b11111111110000111000111111111111;
			13'h137c: data = 32'b11111111110000110000111111111111;
			13'h137d: data = 32'b11111111110000110000111111111111;
			13'h137e: data = 32'b11111111110000110000111111111111;
			13'h137f: data = 32'b10000000000000000000000000000000;

//n x4e
			13'h1380: data = 32'b11111111100000000000001111111111;
			13'h1381: data = 32'b11111111110000000000011111111111;
			13'h1382: data = 32'b11111111110000000000011111111111;
			13'h1383: data = 32'b11111111111000000000011111111111;
			13'h1384: data = 32'b11111111111000000000011111111111;
			13'h1385: data = 32'b11111111111100000000011111111111;
			13'h1386: data = 32'b11111111111100000000011111111111;
			13'h1387: data = 32'b11111111111100000000011111111111;
			13'h1388: data = 32'b11111111111110000000011111111111;
			13'h1389: data = 32'b11111111111110000000011111111111;
			13'h138a: data = 32'b11111111111111000000011111111111;
			13'h138b: data = 32'b11111111111111000000011111111111;
			13'h138c: data = 32'b11111111111111000000011111111111;
			13'h138d: data = 32'b11111111111111100000011111111111;
			13'h138e: data = 32'b11111111111111100000011111111111;
			13'h138f: data = 32'b11111111111111110000011111111111;
			13'h1390: data = 32'b11111111111111110000011111111111;
			13'h1391: data = 32'b11111111111111110000011111111111;
			13'h1392: data = 32'b11111111111111111000011111111111;
			13'h1393: data = 32'b11111111111111111000011111111111;
			13'h1394: data = 32'b11111111111111111100011111111111;
			13'h1395: data = 32'b11111111111111111100011111111111;
			13'h1396: data = 32'b11111111111111111100011111111111;
			13'h1397: data = 32'b11111111111111111110011111111111;
			13'h1398: data = 32'b11111111111111111110011111111111;
			13'h1399: data = 32'b11111111111111111111011111111111;
			13'h139a: data = 32'b11111111111111111111011111111111;
			13'h139b: data = 32'b11111111111111111111011111111111;
			13'h139c: data = 32'b11111111111111111111101111111111;
			13'h139d: data = 32'b11111111111111111111101111111111;
			13'h139e: data = 32'b11111111111111111111111111111111;
			13'h139f: data = 32'b11111111111111111111111111111111;
			13'h13a0: data = 32'b11111111111111111111111111111111;
			13'h13a1: data = 32'b11111111111111111111111111111111;
			13'h13a2: data = 32'b11111111110111111111111111111111;
			13'h13a3: data = 32'b11111111110111111111111111111111;
			13'h13a4: data = 32'b11111111110111111111111111111111;
			13'h13a5: data = 32'b11111111110011111111111111111111;
			13'h13a6: data = 32'b11111111110011111111111111111111;
			13'h13a7: data = 32'b11111111110001111111111111111111;
			13'h13a8: data = 32'b11111111110001111111111111111111;
			13'h13a9: data = 32'b11111111110001111111111111111111;
			13'h13aa: data = 32'b11111111110000111111111111111111;
			13'h13ab: data = 32'b11111111110000111111111111111111;
			13'h13ac: data = 32'b11111111110000011111111111111111;
			13'h13ad: data = 32'b11111111110000011111111111111111;
			13'h13ae: data = 32'b11111111110000001111111111111111;
			13'h13af: data = 32'b11111111110000001111111111111111;
			13'h13b0: data = 32'b11111111110000001111111111111111;
			13'h13b1: data = 32'b11111111110000000111111111111111;
			13'h13b2: data = 32'b11111111110000000111111111111111;
			13'h13b3: data = 32'b11111111110000000011111111111111;
			13'h13b4: data = 32'b11111111110000000011111111111111;
			13'h13b5: data = 32'b11111111110000000011111111111111;
			13'h13b6: data = 32'b11111111110000000001111111111111;
			13'h13b7: data = 32'b11111111110000000001111111111111;
			13'h13b8: data = 32'b11111111110000000000111111111111;
			13'h13b9: data = 32'b11111111110000000000111111111111;
			13'h13ba: data = 32'b11111111110000000000111111111111;
			13'h13bb: data = 32'b11111111110000000000011111111111;
			13'h13bc: data = 32'b11111111110000000000011111111111;
			13'h13bd: data = 32'b11111111110000000000001111111111;
			13'h13be: data = 32'b11111111110000000000001111111111;
			13'h13bf: data = 32'b00000000000000000000000000000000;

//O x4f
			13'h13c0: data = 32'b00000000000000000000000000000000;
			13'h13c1: data = 32'b00000000000000111110000000000000;
			13'h13c2: data = 32'b00000000000011111111100000000000;
			13'h13c3: data = 32'b00000000000111111111110000000000;
			13'h13c4: data = 32'b00000000001111111111111000000000;
			13'h13c5: data = 32'b00000000011111111111111100000000;
			13'h13c6: data = 32'b00000000111111111111111110000000;
			13'h13c7: data = 32'b00000001111111100011111111000000;
			13'h13c8: data = 32'b00000001111111000001111111000000;
			13'h13c9: data = 32'b00000011111110000000111111100000;
			13'h13ca: data = 32'b00000011111100000000011111100000;
			13'h13cb: data = 32'b00000111111100000000011111110000;
			13'h13cc: data = 32'b00000111111000000000001111110000;
			13'h13cd: data = 32'b00000111111000000000001111110000;
			13'h13ce: data = 32'b00001111110000000000001111111000;
			13'h13cf: data = 32'b00001111110000000000000111111000;
			13'h13d0: data = 32'b00001111110000000000000111111000;
			13'h13d1: data = 32'b00011111110000000000000111111000;
			13'h13d2: data = 32'b00011111100000000000000111111100;
			13'h13d3: data = 32'b00011111100000000000000011111100;
			13'h13d4: data = 32'b00011111100000000000000011111100;
			13'h13d5: data = 32'b00011111100000000000000011111100;
			13'h13d6: data = 32'b00011111100000000000000011111100;
			13'h13d7: data = 32'b00111111100000000000000011111100;
			13'h13d8: data = 32'b00111111100000000000000011111110;
			13'h13d9: data = 32'b00111111100000000000000011111110;
			13'h13da: data = 32'b00111111100000000000000011111110;
			13'h13db: data = 32'b00111111100000000000000011111110;
			13'h13dc: data = 32'b00111111100000000000000011111110;
			13'h13dd: data = 32'b00111111100000000000000011111110;
			13'h13de: data = 32'b00111111100000000000000011111110;
			13'h13df: data = 32'b00111111100000000000000011111110;
			13'h13e0: data = 32'b00111111100000000000000011111110;
			13'h13e1: data = 32'b00111111100000000000000011111110;
			13'h13e2: data = 32'b00111111100000000000000011111110;
			13'h13e3: data = 32'b00111111100000000000000011111110;
			13'h13e4: data = 32'b00111111100000000000000011111110;
			13'h13e5: data = 32'b00111111100000000000000011111110;
			13'h13e6: data = 32'b00111111100000000000000011111110;
			13'h13e7: data = 32'b00111111100000000000000011111110;
			13'h13e8: data = 32'b00111111100000000000000011111100;
			13'h13e9: data = 32'b00011111100000000000000011111100;
			13'h13ea: data = 32'b00011111100000000000000011111100;
			13'h13eb: data = 32'b00011111100000000000000011111100;
			13'h13ec: data = 32'b00011111100000000000000011111100;
			13'h13ed: data = 32'b00011111100000000000000111111100;
			13'h13ee: data = 32'b00011111110000000000000111111000;
			13'h13ef: data = 32'b00001111110000000000000111111000;
			13'h13f0: data = 32'b00001111110000000000000111111000;
			13'h13f1: data = 32'b00001111110000000000001111111000;
			13'h13f2: data = 32'b00000111111000000000001111110000;
			13'h13f3: data = 32'b00000111111000000000001111110000;
			13'h13f4: data = 32'b00000111111100000000011111100000;
			13'h13f5: data = 32'b00000011111100000000011111100000;
			13'h13f6: data = 32'b00000011111110000000111111000000;
			13'h13f7: data = 32'b00000001111111000001111111000000;
			13'h13f8: data = 32'b00000001111111111111111110000000;
			13'h13f9: data = 32'b00000000111111111111111110000000;
			13'h13fa: data = 32'b00000000011111111111111100000000;


//P x50
			13'h1400: data = 32'b01111111111111111110000000000000;
			13'h1401: data = 32'b01111111111111111111100000000000;
			13'h1402: data = 32'b01111111111111111111111000000000;
			13'h1403: data = 32'b00111111111111111111111100000000;
			13'h1404: data = 32'b00001111111111111111111110000000;
			13'h1405: data = 32'b00001111111100001111111111000000;
			13'h1406: data = 32'b00000111111100000011111111100000;
			13'h1407: data = 32'b00000111111100000001111111100000;
			13'h1408: data = 32'b00000111111100000000111111110000;
			13'h1409: data = 32'b00000111111100000000011111110000;
			13'h140a: data = 32'b00000111111100000000001111111000;
			13'h140b: data = 32'b00000111111100000000001111111000;
			13'h140c: data = 32'b00000111111100000000001111111000;
			13'h140d: data = 32'b00000111111100000000000111111000;
			13'h140e: data = 32'b00000111111100000000000111111100;
			13'h140f: data = 32'b00000111111100000000000111111100;
			13'h1410: data = 32'b00000111111100000000000111111100;
			13'h1411: data = 32'b00000111111100000000000111111100;
			13'h1412: data = 32'b00000111111100000000000111111100;
			13'h1413: data = 32'b00000111111100000000000111111100;
			13'h1414: data = 32'b00000111111100000000000111111100;
			13'h1415: data = 32'b00000111111100000000000111111100;
			13'h1416: data = 32'b00000111111100000000000111111100;
			13'h1417: data = 32'b00000111111100000000000111111100;
			13'h1418: data = 32'b00000111111100000000000111111000;
			13'h1419: data = 32'b00000111111100000000001111111000;
			13'h141a: data = 32'b00000111111100000000001111111000;
			13'h141b: data = 32'b00000111111100000000001111111000;
			13'h141c: data = 32'b00000111111100000000011111110000;
			13'h141d: data = 32'b00000111111100000000111111110000;
			13'h141e: data = 32'b00000111111100000001111111100000;
			13'h141f: data = 32'b00000111111100001111111111100000;
			13'h1420: data = 32'b00000111111111111111111111000000;
			13'h1421: data = 32'b00000111111111111111111110000000;
			13'h1422: data = 32'b00000111111111111111111100000000;
			13'h1423: data = 32'b00000111111111111111110000000000;
			13'h1424: data = 32'b00000111111111111111000000000000;
			13'h1425: data = 32'b00000111111111000000000000000000;
			13'h1426: data = 32'b00000111111100000000000000000000;
			13'h1427: data = 32'b00000111111100000000000000000000;
			13'h1428: data = 32'b00000111111100000000000000000000;
			13'h1429: data = 32'b00000111111100000000000000000000;
			13'h142a: data = 32'b00000111111100000000000000000000;
			13'h142b: data = 32'b00000111111100000000000000000000;
			13'h142c: data = 32'b00000111111100000000000000000000;
			13'h142d: data = 32'b00000111111100000000000000000000;
			13'h142e: data = 32'b00000111111100000000000000000000;
			13'h142f: data = 32'b00000111111100000000000000000000;
			13'h1430: data = 32'b00000111111100000000000000000000;
			13'h1431: data = 32'b00000111111100000000000000000000;
			13'h1432: data = 32'b00000111111100000000000000000000;
			13'h1433: data = 32'b00000111111100000000000000000000;
			13'h1434: data = 32'b00000111111100000000000000000000;
			13'h1435: data = 32'b00000111111100000000000000000000;
			13'h1436: data = 32'b00000111111100000000000000000000;
			13'h1437: data = 32'b00000111111100000000000000000000;
			13'h1438: data = 32'b00000111111100000000000000000000;
			13'h1439: data = 32'b00000111111100000000000000000000;
			13'h143a: data = 32'b00000111111100000000000000000000;
			13'h143b: data = 32'b00001111111110000000000000000000;
			13'h143c: data = 32'b01111111111111110000000000000000;
			13'h143d: data = 32'b11111111111111110000000000000000;
			13'h143e: data = 32'b11111111111111110000000000000000;
			13'h143f: data = 32'b11111111111111110000000000000000;
			13'h13fb: data = 32'b00000000001111111111111000000000;
			13'h13fc: data = 32'b00000000000111111111110000000000;
			13'h13fd: data = 32'b00000000000011111111000000000000;
			13'h13fe: data = 32'b00000000000000011100000000000000;
			13'h13ff: data = 32'b00000000000000000000000000000000;

//p x51
			13'h1440: data = 32'b00000000000001111110000000000000;
			13'h1441: data = 32'b00000000000111111111100000000000;
			13'h1442: data = 32'b00000000001111111111110000000000;
			13'h1443: data = 32'b00000000011111111111111000000000;
			13'h1444: data = 32'b00000000111111111111111100000000;
			13'h1445: data = 32'b00000001111111000111111100000000;
			13'h1446: data = 32'b00000001111110000001111110000000;
			13'h1447: data = 32'b00000011111100000001111110000000;
			13'h1448: data = 32'b00000011111100000000111111000000;
			13'h1449: data = 32'b00000111111000000000011111000000;
			13'h144a: data = 32'b00000111111000000000011111100000;
			13'h144b: data = 32'b00000111110000000000011111100000;
			13'h144c: data = 32'b00001111110000000000001111100000;
			13'h144d: data = 32'b00001111110000000000001111110000;
			13'h144e: data = 32'b00001111110000000000001111110000;
			13'h144f: data = 32'b00001111100000000000001111110000;
			13'h1450: data = 32'b00011111100000000000001111110000;
			13'h1451: data = 32'b00011111100000000000000111110000;
			13'h1452: data = 32'b00011111100000000000000111111000;
			13'h1453: data = 32'b00011111100000000000000111111000;
			13'h1454: data = 32'b00011111100000000000000111111000;
			13'h1455: data = 32'b00011111100000000000000111111000;
			13'h1456: data = 32'b00011111100000000000000111111000;
			13'h1457: data = 32'b00011111100000000000000111111000;
			13'h1458: data = 32'b00011111100000000000000111111000;
			13'h1459: data = 32'b00011111100000000000000111111000;
			13'h145a: data = 32'b00011111100000000000000111111000;
			13'h145b: data = 32'b00011111100000000000000111111000;
			13'h145c: data = 32'b00011111100000000000000111111000;
			13'h145d: data = 32'b00011111100000000000000111111000;
			13'h145e: data = 32'b00011111100000000000000111111000;
			13'h145f: data = 32'b00011111100000000000000111111000;
			13'h1460: data = 32'b00011111100000000000000111111000;
			13'h1461: data = 32'b00011111100000000000000111111000;
			13'h1462: data = 32'b00011111100000000000000111111000;
			13'h1463: data = 32'b00011111100000000000000111110000;
			13'h1464: data = 32'b00001111100000000000001111110000;
			13'h1465: data = 32'b00001111110000000000001111110000;
			13'h1466: data = 32'b00001111110000000000001111110000;
			13'h1467: data = 32'b00001111110000000000001111100000;
			13'h1468: data = 32'b00000111110000000000001111100000;
			13'h1469: data = 32'b00000111111000000000011111100000;
			13'h146a: data = 32'b00000111111000000000011111100000;
			13'h146b: data = 32'b00000011111000000000111111000000;
			13'h146c: data = 32'b00000011111100000000111111000000;
			13'h146d: data = 32'b00000001111110000001111110000000;
			13'h146e: data = 32'b00000001111111000011111110000000;
			13'h146f: data = 32'b00000000111111111111111100000000;
			13'h1470: data = 32'b00000000011111111111111000000000;
			13'h1471: data = 32'b00000000001111111111110000000000;
			13'h1472: data = 32'b00000000001111111111100000000000;
			13'h1473: data = 32'b00000000000011111111000000000000;
			13'h1474: data = 32'b00000000000011111111000000000000;
			13'h1475: data = 32'b00000000000001111111000000000000;
			13'h1476: data = 32'b00000000000001111111100000000000;
			13'h1477: data = 32'b00000000000000111111110000000000;
			13'h1478: data = 32'b00000000000000111111110000000000;
			13'h1479: data = 32'b00000000000000011111111000000000;
			13'h147a: data = 32'b00000000000000011111111100000000;
			13'h147b: data = 32'b00000000000000001111111111000000;
			13'h147c: data = 32'b00000000000000000111111111111000;
			13'h147d: data = 32'b00000000000000000011111111111100;
			13'h147e: data = 32'b00000000000000000000111111111100;
			13'h147f: data = 32'b00000000000000000000001111111100;

//R x52 R
			13'h1480: data = 32'b00000000000000000000000000000000;
			13'h1481: data = 32'b01111111111111111111100000000000;
			13'h1482: data = 32'b01111111111111111111111000000000;
			13'h1483: data = 32'b01111111111111111111111100000000;
			13'h1484: data = 32'b01111111111111111111111110000000;
			13'h1485: data = 32'b01111111111111111111111111000000;
			13'h1486: data = 32'b01111111111111111111111111000000;
			13'h1487: data = 32'b01111111111111111111111111100000;
			13'h1488: data = 32'b01111111111111111111111111100000;
			13'h1489: data = 32'b01111111111111111111111111110000;
			13'h148a: data = 32'b01111111111111111111111111110000;
			13'h148b: data = 32'b01111111111111111111111111110000;
			13'h148c: data = 32'b01111111000000000001111111110000;
			13'h148d: data = 32'b01111111100000000000111111110000;
			13'h148e: data = 32'b01111111100000000000111111111000;
			13'h148f: data = 32'b01111111100000000000011111111000;
			13'h1490: data = 32'b01111111100000000000011111111000;
			13'h1491: data = 32'b01111111100000000000011111111000;
			13'h1492: data = 32'b01111111100000000000011111111000;
			13'h1493: data = 32'b01111111100000000000011111111000;
			13'h1494: data = 32'b01111111100000000000011111111000;
			13'h1495: data = 32'b01111111100000000000011111111000;
			13'h1496: data = 32'b01111111100000000000011111111000;
			13'h1497: data = 32'b01111111100000000000011111110000;
			13'h1498: data = 32'b01111111100000000000111111110000;
			13'h1499: data = 32'b01111111100000000000111111110000;
			13'h149a: data = 32'b01111111000000000011111111110000;
			13'h149b: data = 32'b01111111111111111111111111110000;
			13'h149c: data = 32'b01111111111111111111111111100000;
			13'h149d: data = 32'b01111111111111111111111111100000;
			13'h149e: data = 32'b01111111111111111111111111000000;
			13'h149f: data = 32'b01111111111111111111111111000000;
			13'h14a0: data = 32'b01111111111111111111111110000000;
			13'h14a1: data = 32'b01111111111111111111111100000000;
			13'h14a2: data = 32'b01111111111111111111111000000000;
			13'h14a3: data = 32'b01111111111111111111100000000000;
			13'h14a4: data = 32'b01111111111111111111100000000000;
			13'h14a5: data = 32'b01111111000011111111110000000000;
			13'h14a6: data = 32'b01111111100001111111110000000000;
			13'h14a7: data = 32'b01111111100000111111111000000000;
			13'h14a8: data = 32'b01111111100000011111111100000000;
			13'h14a9: data = 32'b01111111100000011111111100000000;
			13'h14aa: data = 32'b01111111100000011111111110000000;
			13'h14ab: data = 32'b01111111100000001111111110000000;
			13'h14ac: data = 32'b01111111100000001111111110000000;
			13'h14ad: data = 32'b01111111100000000111111111000000;
			13'h14ae: data = 32'b01111111100000000111111111000000;
			13'h14af: data = 32'b01111111100000000111111111000000;
			13'h14b0: data = 32'b01111111100000000011111111100000;
			13'h14b1: data = 32'b01111111100000000011111111100000;
			13'h14b2: data = 32'b01111111100000000011111111100000;
			13'h14b3: data = 32'b01111111100000000001111111110000;
			13'h14b4: data = 32'b01111111100000000001111111110000;
			13'h14b5: data = 32'b01111111100000000000111111110000;
			13'h14b6: data = 32'b01111111100000000000111111111000;
			13'h14b7: data = 32'b01111111100000000000111111111000;
			13'h14b8: data = 32'b01111111100000000000011111111000;
			13'h14b9: data = 32'b01111111100000000000011111111100;
			13'h14ba: data = 32'b01111111100000000000011111111100;
			13'h14bb: data = 32'b01111111100000000000001111111100;
			13'h14bc: data = 32'b01111111100000000000001111111110;
			13'h14bd: data = 32'b01111111100000000000001111111110;
			13'h14be: data = 32'b01111111100000000000000111111110;
			13'h14bf: data = 32'b00000000000000000000000000000000;

//S x53
			13'h14c0: data = 32'b00000000000000011100000000000000;
			13'h14c1: data = 32'b00000000000111111111110000000000;
			13'h14c2: data = 32'b00000000001111111111111100000000;
			13'h14c3: data = 32'b00000000011111111111111111000000;
			13'h14c4: data = 32'b00000000111111111111111111100000;
			13'h14c5: data = 32'b00000001111111111111111111110000;
			13'h14c6: data = 32'b00000011111111111111111111111000;
			13'h14c7: data = 32'b00000011111111111111111111111000;
			13'h14c8: data = 32'b00000111111111111111111111111000;
			13'h14c9: data = 32'b00000111111111111111111111111000;
			13'h14ca: data = 32'b00001111111111111111111111111000;
			13'h14cb: data = 32'b00001111111111111111111111111000;
			13'h14cc: data = 32'b00001111111111111111111111111000;
			13'h14cd: data = 32'b00001111111111111111111111110000;
			13'h14ce: data = 32'b00011111111111111111111111110000;
			13'h14cf: data = 32'b00011111111111111111111111110000;
			13'h14d0: data = 32'b00011111111111100000111111110000;
			13'h14d1: data = 32'b00011111111111000000001111110000;
			13'h14d2: data = 32'b00011111111111000000000011100000;
			13'h14d3: data = 32'b00011111111111100000000001100000;
			13'h14d4: data = 32'b00011111111111100000000000100000;
			13'h14d5: data = 32'b00011111111111111000000000000000;
			13'h14d6: data = 32'b00011111111111111110000000000000;
			13'h14d7: data = 32'b00011111111111111111100000000000;
			13'h14d8: data = 32'b00011111111111111111111000000000;
			13'h14d9: data = 32'b00011111111111111111111100000000;
			13'h14da: data = 32'b00001111111111111111111111000000;
			13'h14db: data = 32'b00001111111111111111111111100000;
			13'h14dc: data = 32'b00001111111111111111111111100000;
			13'h14dd: data = 32'b00001111111111111111111111110000;
			13'h14de: data = 32'b00000111111111111111111111111000;
			13'h14df: data = 32'b00000111111111111111111111111000;
			13'h14e0: data = 32'b00000011111111111111111111111000;
			13'h14e1: data = 32'b00000011111111111111111111111100;
			13'h14e2: data = 32'b00000001111111111111111111111100;
			13'h14e3: data = 32'b00000000111111111111111111111100;
			13'h14e4: data = 32'b00000000011111111111111111111110;
			13'h14e5: data = 32'b00000000001111111111111111111110;
			13'h14e6: data = 32'b00000000000111111111111111111110;
			13'h14e7: data = 32'b00000000000001111111111111111110;
			13'h14e8: data = 32'b00000000000000011111111111111110;
			13'h14e9: data = 32'b00001100000000000111111111111110;
			13'h14ea: data = 32'b00001110000000000001111111111110;
			13'h14eb: data = 32'b00001111000000000001111111111110;
			13'h14ec: data = 32'b00001111100000000000111111111110;
			13'h14ed: data = 32'b00001111110000000000111111111110;
			13'h14ee: data = 32'b00001111111000000001111111111110;
			13'h14ef: data = 32'b00011111111110000001111111111110;
			13'h14f0: data = 32'b00011111111111111111111111111110;
			13'h14f1: data = 32'b00011111111111111111111111111110;
			13'h14f2: data = 32'b00011111111111111111111111111100;
			13'h14f3: data = 32'b00011111111111111111111111111100;
			13'h14f4: data = 32'b00011111111111111111111111111100;
			13'h14f5: data = 32'b00111111111111111111111111111100;
			13'h14f6: data = 32'b00111111111111111111111111111000;
			13'h14f7: data = 32'b00111111111111111111111111111000;
			13'h14f8: data = 32'b00011111111111111111111111110000;
			13'h14f9: data = 32'b00001111111111111111111111110000;
			13'h14fa: data = 32'b00000111111111111111111111100000;
			13'h14fb: data = 32'b00000011111111111111111111000000;
			13'h14fc: data = 32'b00000001111111111111111110000000;
			13'h14fd: data = 32'b00000000011111111111111100000000;
			13'h14fe: data = 32'b00000000000111111111110000000000;
			13'h14ff: data = 32'b00000000000000111110000000000000;


//T x54
			13'h1500: data = 32'b00000000000000000000000000000000;
			13'h1501: data = 32'b01111111111111111111111111111110;
			13'h1502: data = 32'b01111111111111111111111111111110;
			13'h1503: data = 32'b01111111111111111111111111111110;
			13'h1504: data = 32'b01111111111111111111111111111110;
			13'h1505: data = 32'b01111111111111111111111111111110;
			13'h1506: data = 32'b01111111111111111111111111111110;
			13'h1507: data = 32'b01111111111111111111111111111110;
			13'h1508: data = 32'b01111111111111111111111111111110;
			13'h1509: data = 32'b01111111111111111111111111111110;
			13'h150a: data = 32'b01111111111111111111111111111110;
			13'h150b: data = 32'b01111111111111111111111111111110;
			13'h150c: data = 32'b01111111111111111111111111111110;
			13'h150d: data = 32'b01111111111111111111111111111110;
			13'h150e: data = 32'b01111111111111111111111111111110;
			13'h150f: data = 32'b01111111111111111111111111111110;
			13'h1510: data = 32'b00000000000111111111110000000000;
			13'h1511: data = 32'b00000000000111111111110000000000;
			13'h1512: data = 32'b00000000000111111111110000000000;
			13'h1513: data = 32'b00000000000111111111110000000000;
			13'h1514: data = 32'b00000000000111111111110000000000;
			13'h1515: data = 32'b00000000000111111111110000000000;
			13'h1516: data = 32'b00000000000111111111110000000000;
			13'h1517: data = 32'b00000000000111111111110000000000;
			13'h1518: data = 32'b00000000000111111111110000000000;
			13'h1519: data = 32'b00000000000111111111110000000000;
			13'h151a: data = 32'b00000000000111111111110000000000;
			13'h151b: data = 32'b00000000000111111111110000000000;
			13'h151c: data = 32'b00000000000111111111110000000000;
			13'h151d: data = 32'b00000000000111111111110000000000;
			13'h151e: data = 32'b00000000000111111111110000000000;
			13'h151f: data = 32'b00000000000111111111110000000000;
			13'h1520: data = 32'b00000000000111111111110000000000;
			13'h1521: data = 32'b00000000000111111111110000000000;
			13'h1522: data = 32'b00000000000111111111110000000000;
			13'h1523: data = 32'b00000000000111111111110000000000;
			13'h1524: data = 32'b00000000000111111111110000000000;
			13'h1525: data = 32'b00000000000111111111110000000000;
			13'h1526: data = 32'b00000000000111111111110000000000;
			13'h1527: data = 32'b00000000000111111111110000000000;
			13'h1528: data = 32'b00000000000111111111110000000000;
			13'h1529: data = 32'b00000000000111111111110000000000;
			13'h152a: data = 32'b00000000000111111111110000000000;
			13'h152b: data = 32'b00000000000111111111110000000000;
			13'h152c: data = 32'b00000000000111111111110000000000;
			13'h152d: data = 32'b00000000000111111111110000000000;
			13'h152e: data = 32'b00000000000111111111110000000000;
			13'h152f: data = 32'b00000000000111111111110000000000;
			13'h1530: data = 32'b00000000000111111111110000000000;
			13'h1531: data = 32'b00000000000111111111110000000000;
			13'h1532: data = 32'b00000000000111111111110000000000;
			13'h1533: data = 32'b00000000000111111111110000000000;
			13'h1534: data = 32'b00000000000111111111110000000000;
			13'h1535: data = 32'b00000000000111111111110000000000;
			13'h1536: data = 32'b00000000000111111111110000000000;
			13'h1537: data = 32'b00000000000111111111110000000000;
			13'h1538: data = 32'b00000000000111111111110000000000;
			13'h1539: data = 32'b00000000000111111111110000000000;
			13'h153a: data = 32'b00000000000111111111110000000000;
			13'h153b: data = 32'b00000000000111111111110000000000;
			13'h153c: data = 32'b00000000000111111111110000000000;
			13'h153d: data = 32'b00000000000111111111110000000000;
			13'h153e: data = 32'b00000000000111111111110000000000;
			13'h153f: data = 32'b00000000000000000000000000000000;


// U x55
			13'h1540: data = 32'b00000000000000000000000000000000;
			13'h1541: data = 32'b00000000000000000000000000000000;
			13'h1542: data = 32'b00111111111111100000111111111111;
			13'h1543: data = 32'b00111111111111100000111111111111;
			13'h1544: data = 32'b00111111111111100000111111111111;
			13'h1545: data = 32'b00111111111111100000111111111111;
			13'h1546: data = 32'b00111111111111100000011111111111;
			13'h1547: data = 32'b00000111111100000000000111111000;
			13'h1548: data = 32'b00000111111100000000000011110000;
			13'h1549: data = 32'b00000111111000000000000011110000;
			13'h154a: data = 32'b00000111111000000000000011110000;
			13'h154b: data = 32'b00000111111000000000000011110000;
			13'h154c: data = 32'b00000111111000000000000011110000;
			13'h154d: data = 32'b00000111111000000000000011110000;
			13'h154e: data = 32'b00000111111000000000000011110000;
			13'h154f: data = 32'b00000111111000000000000011110000;
			13'h1550: data = 32'b00000111111000000000000011110000;
			13'h1551: data = 32'b00000111111000000000000011110000;
			13'h1552: data = 32'b00000111111000000000000011110000;
			13'h1553: data = 32'b00000111111000000000000011110000;
			13'h1554: data = 32'b00000111111000000000000011110000;
			13'h1555: data = 32'b00000111111000000000000011110000;
			13'h1556: data = 32'b00000111111000000000000011110000;
			13'h1557: data = 32'b00000111111000000000000011110000;
			13'h1558: data = 32'b00000111111000000000000011110000;
			13'h1559: data = 32'b00000111111000000000000011110000;
			13'h155a: data = 32'b00000111111000000000000011110000;
			13'h155b: data = 32'b00000111111000000000000011110000;
			13'h155c: data = 32'b00000111111000000000000011110000;
			13'h155d: data = 32'b00000111111000000000000011110000;
			13'h155e: data = 32'b00000111111000000000000011110000;
			13'h155f: data = 32'b00000111111000000000000011110000;
			13'h1560: data = 32'b00000111111000000000000011110000;
			13'h1561: data = 32'b00000111111000000000000011110000;
			13'h1562: data = 32'b00000111111000000000000011110000;
			13'h1563: data = 32'b00000111111000000000000011110000;
			13'h1564: data = 32'b00000111111000000000000011110000;
			13'h1565: data = 32'b00000111111000000000000011110000;
			13'h1566: data = 32'b00000111111000000000000011110000;
			13'h1567: data = 32'b00000111111000000000000011110000;
			13'h1568: data = 32'b00000111111000000000000011110000;
			13'h1569: data = 32'b00000111111000000000000011110000;
			13'h156a: data = 32'b00000111111000000000000011110000;
			13'h156b: data = 32'b00000111111000000000000011110000;
			13'h156c: data = 32'b00000111111000000000000011110000;
			13'h156d: data = 32'b00000111111100000000000011110000;
			13'h156e: data = 32'b00000011111100000000000011110000;
			13'h156f: data = 32'b00000011111100000000000011100000;
			13'h1570: data = 32'b00000011111100000000000111100000;
			13'h1571: data = 32'b00000011111100000000000111100000;
			13'h1572: data = 32'b00000011111100000000000111100000;
			13'h1573: data = 32'b00000011111110000000000111100000;
			13'h1574: data = 32'b00000001111110000000001111000000;
			13'h1575: data = 32'b00000001111111000000011111000000;
			13'h1576: data = 32'b00000001111111100000111111000000;
			13'h1577: data = 32'b00000000111111111111111110000000;
			13'h1578: data = 32'b00000000111111111111111110000000;
			13'h1579: data = 32'b00000000011111111111111100000000;
			13'h157a: data = 32'b00000000001111111111111000000000;
			13'h157b: data = 32'b00000000000111111111110000000000;
			13'h157c: data = 32'b00000000000011111111100000000000;
			13'h157d: data = 32'b00000000000000111110000000000000;
			13'h157e: data = 32'b00000000000000000000000000000000;
			13'h157f: data = 32'b00000000000000000000000000000000;



//Y x59
			13'h1640: data = 32'b00000000000000000000000000000000;
			13'h1641: data = 32'b00000000000000000000000000000001;
			13'h1642: data = 32'b11111111111000000000011111111111;
			13'h1643: data = 32'b11111111111000000000011111111111;
			13'h1644: data = 32'b01111111111000000000111111111110;
			13'h1645: data = 32'b01111111111100000000111111111110;
			13'h1646: data = 32'b01111111111100000000111111111110;
			13'h1647: data = 32'b00111111111100000000111111111100;
			13'h1648: data = 32'b00111111111110000001111111111100;
			13'h1649: data = 32'b00111111111110000001111111111100;
			13'h164a: data = 32'b00111111111110000001111111111000;
			13'h164b: data = 32'b00011111111110000011111111111000;
			13'h164c: data = 32'b00011111111111000011111111111000;
			13'h164d: data = 32'b00011111111111000011111111110000;
			13'h164e: data = 32'b00001111111111000011111111110000;
			13'h164f: data = 32'b00001111111111100111111111110000;
			13'h1650: data = 32'b00001111111111100111111111110000;
			13'h1651: data = 32'b00000111111111100111111111100000;
			13'h1652: data = 32'b00000111111111101111111111100000;
			13'h1653: data = 32'b00000111111111111111111111100000;
			13'h1654: data = 32'b00000011111111111111111111000000;
			13'h1655: data = 32'b00000011111111111111111111000000;
			13'h1656: data = 32'b00000011111111111111111111000000;
			13'h1657: data = 32'b00000011111111111111111110000000;
			13'h1658: data = 32'b00000001111111111111111110000000;
			13'h1659: data = 32'b00000001111111111111111110000000;
			13'h165a: data = 32'b00000001111111111111111100000000;
			13'h165b: data = 32'b00000000111111111111111100000000;
			13'h165c: data = 32'b00000000111111111111111100000000;
			13'h165d: data = 32'b00000000111111111111111000000000;
			13'h165e: data = 32'b00000000011111111111111000000000;
			13'h165f: data = 32'b00000000011111111111111000000000;
			13'h1660: data = 32'b00000000011111111111110000000000;
			13'h1661: data = 32'b00000000001111111111110000000000;
			13'h1662: data = 32'b00000000001111111111110000000000;
			13'h1663: data = 32'b00000000001111111111110000000000;
			13'h1664: data = 32'b00000000001111111111100000000000;
			13'h1665: data = 32'b00000000000111111111100000000000;
			13'h1666: data = 32'b00000000000111111111100000000000;
			13'h1667: data = 32'b00000000000111111111100000000000;
			13'h1668: data = 32'b00000000000111111111100000000000;
			13'h1669: data = 32'b00000000000111111111100000000000;
			13'h166a: data = 32'b00000000000111111111100000000000;
			13'h166b: data = 32'b00000000000111111111100000000000;
			13'h166c: data = 32'b00000000000111111111100000000000;
			13'h166d: data = 32'b00000000000111111111100000000000;
			13'h166e: data = 32'b00000000000111111111100000000000;
			13'h166f: data = 32'b00000000000111111111100000000000;
			13'h1670: data = 32'b00000000000111111111100000000000;
			13'h1671: data = 32'b00000000000111111111100000000000;
			13'h1672: data = 32'b00000000000111111111100000000000;
			13'h1673: data = 32'b00000000000111111111100000000000;
			13'h1674: data = 32'b00000000000111111111100000000000;
			13'h1675: data = 32'b00000000000111111111100000000000;
			13'h1676: data = 32'b00000000000111111111100000000000;
			13'h1677: data = 32'b00000000000111111111100000000000;
			13'h1678: data = 32'b00000000000111111111100000000000;
			13'h1679: data = 32'b00000000000111111111100000000000;
			13'h167a: data = 32'b00000000000111111111100000000000;
			13'h167b: data = 32'b00000000000111111111100000000000;
			13'h167c: data = 32'b00000000000111111111100000000000;
			13'h167d: data = 32'b00000000000111111111100000000000;
			13'h167e: data = 32'b00000000000000000000000000000000;
			13'h167f: data = 32'b00000000000000000000000000000000;
			default: data = 32'b00000000000000000000000000000000;

			  endcase  
							 
endmodule      
	       
	